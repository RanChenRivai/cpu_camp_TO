magic
tech sky130A
magscale 1 2
timestamp 1663424475
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 322934 700748 322940 700800
rect 322992 700788 322998 700800
rect 348786 700788 348792 700800
rect 322992 700760 348792 700788
rect 322992 700748 322998 700760
rect 348786 700748 348792 700760
rect 348844 700748 348850 700800
rect 283834 700680 283840 700732
rect 283892 700720 283898 700732
rect 328454 700720 328460 700732
rect 283892 700692 328460 700720
rect 283892 700680 283898 700692
rect 328454 700680 328460 700692
rect 328512 700680 328518 700732
rect 318794 700612 318800 700664
rect 318852 700652 318858 700664
rect 413646 700652 413652 700664
rect 318852 700624 413652 700652
rect 318852 700612 318858 700624
rect 413646 700612 413652 700624
rect 413704 700612 413710 700664
rect 218974 700544 218980 700596
rect 219032 700584 219038 700596
rect 332594 700584 332600 700596
rect 219032 700556 332600 700584
rect 219032 700544 219038 700556
rect 332594 700544 332600 700556
rect 332652 700544 332658 700596
rect 154114 700476 154120 700528
rect 154172 700516 154178 700528
rect 338114 700516 338120 700528
rect 154172 700488 338120 700516
rect 154172 700476 154178 700488
rect 338114 700476 338120 700488
rect 338172 700476 338178 700528
rect 89162 700408 89168 700460
rect 89220 700448 89226 700460
rect 342254 700448 342260 700460
rect 89220 700420 342260 700448
rect 89220 700408 89226 700420
rect 342254 700408 342260 700420
rect 342312 700408 342318 700460
rect 24302 700340 24308 700392
rect 24360 700380 24366 700392
rect 346394 700380 346400 700392
rect 24360 700352 346400 700380
rect 24360 700340 24366 700352
rect 346394 700340 346400 700352
rect 346452 700340 346458 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 345014 700312 345020 700324
rect 8168 700284 345020 700312
rect 8168 700272 8174 700284
rect 345014 700272 345020 700284
rect 345072 700272 345078 700324
rect 413278 700272 413284 700324
rect 413336 700312 413342 700324
rect 559650 700312 559656 700324
rect 413336 700284 559656 700312
rect 413336 700272 413342 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 300118 700000 300124 700052
rect 300176 700040 300182 700052
rect 301498 700040 301504 700052
rect 300176 700012 301504 700040
rect 300176 700000 300182 700012
rect 301498 700000 301504 700012
rect 301556 700000 301562 700052
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106918 699700 106924 699712
rect 105504 699672 106924 699700
rect 105504 699660 105510 699672
rect 106918 699660 106924 699672
rect 106976 699660 106982 699712
rect 428458 699660 428464 699712
rect 428516 699700 428522 699712
rect 429838 699700 429844 699712
rect 428516 699672 429844 699700
rect 428516 699660 428522 699672
rect 429838 699660 429844 699672
rect 429896 699660 429902 699712
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 303614 696940 303620 696992
rect 303672 696980 303678 696992
rect 580166 696980 580172 696992
rect 303672 696952 580172 696980
rect 303672 696940 303678 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 304994 683136 305000 683188
rect 305052 683176 305058 683188
rect 580166 683176 580172 683188
rect 305052 683148 580172 683176
rect 305052 683136 305058 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 302234 670760 302240 670812
rect 302292 670800 302298 670812
rect 580166 670800 580172 670812
rect 302292 670772 580172 670800
rect 302292 670760 302298 670772
rect 580166 670760 580172 670772
rect 580224 670760 580230 670812
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 351914 670732 351920 670744
rect 3568 670704 351920 670732
rect 3568 670692 3574 670704
rect 351914 670692 351920 670704
rect 351972 670692 351978 670744
rect 3510 656888 3516 656940
rect 3568 656928 3574 656940
rect 350534 656928 350540 656940
rect 3568 656900 350540 656928
rect 3568 656888 3574 656900
rect 350534 656888 350540 656900
rect 350592 656888 350598 656940
rect 298094 643084 298100 643136
rect 298152 643124 298158 643136
rect 580166 643124 580172 643136
rect 298152 643096 580172 643124
rect 298152 643084 298158 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 299474 630640 299480 630692
rect 299532 630680 299538 630692
rect 580166 630680 580172 630692
rect 299532 630652 580172 630680
rect 299532 630640 299538 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3326 618264 3332 618316
rect 3384 618304 3390 618316
rect 356054 618304 356060 618316
rect 3384 618276 356060 618304
rect 3384 618264 3390 618276
rect 356054 618264 356060 618276
rect 356112 618264 356118 618316
rect 296714 616836 296720 616888
rect 296772 616876 296778 616888
rect 580166 616876 580172 616888
rect 296772 616848 580172 616876
rect 296772 616836 296778 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3326 605820 3332 605872
rect 3384 605860 3390 605872
rect 354674 605860 354680 605872
rect 3384 605832 354680 605860
rect 3384 605820 3390 605832
rect 354674 605820 354680 605832
rect 354732 605820 354738 605872
rect 293954 590656 293960 590708
rect 294012 590696 294018 590708
rect 579798 590696 579804 590708
rect 294012 590668 579804 590696
rect 294012 590656 294018 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 295334 576852 295340 576904
rect 295392 576892 295398 576904
rect 580166 576892 580172 576904
rect 295392 576864 580172 576892
rect 295392 576852 295398 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3050 565836 3056 565888
rect 3108 565876 3114 565888
rect 361574 565876 361580 565888
rect 3108 565848 361580 565876
rect 3108 565836 3114 565848
rect 361574 565836 361580 565848
rect 361632 565836 361638 565888
rect 292574 563048 292580 563100
rect 292632 563088 292638 563100
rect 579798 563088 579804 563100
rect 292632 563060 579804 563088
rect 292632 563048 292638 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 358814 553432 358820 553444
rect 3384 553404 358820 553432
rect 3384 553392 3390 553404
rect 358814 553392 358820 553404
rect 358872 553392 358878 553444
rect 288434 536800 288440 536852
rect 288492 536840 288498 536852
rect 580166 536840 580172 536852
rect 288492 536812 580172 536840
rect 288492 536800 288498 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 291194 524424 291200 524476
rect 291252 524464 291258 524476
rect 580166 524464 580172 524476
rect 291252 524436 580172 524464
rect 291252 524424 291258 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3326 514768 3332 514820
rect 3384 514808 3390 514820
rect 365714 514808 365720 514820
rect 3384 514780 365720 514808
rect 3384 514768 3390 514780
rect 365714 514768 365720 514780
rect 365772 514768 365778 514820
rect 287054 510620 287060 510672
rect 287112 510660 287118 510672
rect 580166 510660 580172 510672
rect 287112 510632 580172 510660
rect 287112 510620 287118 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 320174 502936 320180 502988
rect 320232 502976 320238 502988
rect 364334 502976 364340 502988
rect 320232 502948 364340 502976
rect 320232 502936 320238 502948
rect 364334 502936 364340 502948
rect 364392 502936 364398 502988
rect 3234 500964 3240 501016
rect 3292 501004 3298 501016
rect 364334 501004 364340 501016
rect 3292 500976 364340 501004
rect 3292 500964 3298 500976
rect 364334 500964 364340 500976
rect 364392 500964 364398 501016
rect 284294 484372 284300 484424
rect 284352 484412 284358 484424
rect 580166 484412 580172 484424
rect 284352 484384 580172 484412
rect 284352 484372 284358 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 40034 473968 40040 474020
rect 40092 474008 40098 474020
rect 344094 474008 344100 474020
rect 40092 473980 344100 474008
rect 40092 473968 40098 473980
rect 344094 473968 344100 473980
rect 344152 473968 344158 474020
rect 311250 472608 311256 472660
rect 311308 472648 311314 472660
rect 494054 472648 494060 472660
rect 311308 472620 494060 472648
rect 311308 472608 311314 472620
rect 494054 472608 494060 472620
rect 494112 472608 494118 472660
rect 286226 470568 286232 470620
rect 286284 470608 286290 470620
rect 579982 470608 579988 470620
rect 286284 470580 579988 470608
rect 286284 470568 286290 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 106918 469820 106924 469872
rect 106976 469860 106982 469872
rect 339494 469860 339500 469872
rect 106976 469832 339500 469860
rect 106976 469820 106982 469832
rect 339494 469820 339500 469832
rect 339552 469820 339558 469872
rect 169754 468460 169760 468512
rect 169812 468500 169818 468512
rect 334710 468500 334716 468512
rect 169812 468472 334716 468500
rect 169812 468460 169818 468472
rect 334710 468460 334716 468472
rect 334768 468460 334774 468512
rect 234614 467100 234620 467152
rect 234672 467140 234678 467152
rect 330018 467140 330024 467152
rect 234672 467112 330024 467140
rect 234672 467100 234678 467112
rect 330018 467100 330024 467112
rect 330076 467100 330082 467152
rect 301498 465672 301504 465724
rect 301556 465712 301562 465724
rect 325694 465712 325700 465724
rect 301556 465684 325700 465712
rect 301556 465672 301562 465684
rect 325694 465672 325700 465684
rect 325752 465672 325758 465724
rect 316034 464312 316040 464364
rect 316092 464352 316098 464364
rect 428458 464352 428464 464364
rect 316092 464324 428464 464352
rect 316092 464312 316098 464324
rect 428458 464312 428464 464324
rect 428516 464312 428522 464364
rect 277210 464040 277216 464092
rect 277268 464080 277274 464092
rect 435358 464080 435364 464092
rect 277268 464052 435364 464080
rect 277268 464040 277274 464052
rect 435358 464040 435364 464052
rect 435416 464040 435422 464092
rect 215938 463972 215944 464024
rect 215996 464012 216002 464024
rect 380066 464012 380072 464024
rect 215996 463984 380072 464012
rect 215996 463972 216002 463984
rect 380066 463972 380072 463984
rect 380124 463972 380130 464024
rect 220078 463904 220084 463956
rect 220136 463944 220142 463956
rect 387886 463944 387892 463956
rect 220136 463916 387892 463944
rect 220136 463904 220142 463916
rect 387886 463904 387892 463916
rect 387944 463904 387950 463956
rect 217318 463836 217324 463888
rect 217376 463876 217382 463888
rect 392578 463876 392584 463888
rect 217376 463848 392584 463876
rect 217376 463836 217382 463848
rect 392578 463836 392584 463848
rect 392636 463836 392642 463888
rect 280706 463768 280712 463820
rect 280764 463808 280770 463820
rect 457438 463808 457444 463820
rect 280764 463780 457444 463808
rect 280764 463768 280770 463780
rect 457438 463768 457444 463780
rect 457496 463768 457502 463820
rect 13078 463700 13084 463752
rect 13136 463740 13142 463752
rect 378502 463740 378508 463752
rect 13136 463712 378508 463740
rect 13136 463700 13142 463712
rect 378502 463700 378508 463712
rect 378560 463700 378566 463752
rect 235350 462816 235356 462868
rect 235408 462856 235414 462868
rect 375466 462856 375472 462868
rect 235408 462828 375472 462856
rect 235408 462816 235414 462828
rect 375466 462816 375472 462828
rect 375524 462816 375530 462868
rect 264882 462748 264888 462800
rect 264940 462788 264946 462800
rect 422938 462788 422944 462800
rect 264940 462760 422944 462788
rect 264940 462748 264946 462760
rect 422938 462748 422944 462760
rect 422996 462748 423002 462800
rect 221458 462680 221464 462732
rect 221516 462720 221522 462732
rect 383286 462720 383292 462732
rect 221516 462692 383292 462720
rect 221516 462680 221522 462692
rect 383286 462680 383292 462692
rect 383344 462680 383350 462732
rect 260374 462612 260380 462664
rect 260432 462652 260438 462664
rect 421558 462652 421564 462664
rect 260432 462624 421564 462652
rect 260432 462612 260438 462624
rect 421558 462612 421564 462624
rect 421616 462612 421622 462664
rect 279142 462544 279148 462596
rect 279200 462584 279206 462596
rect 454678 462584 454684 462596
rect 279200 462556 454684 462584
rect 279200 462544 279206 462556
rect 454678 462544 454684 462556
rect 454736 462544 454742 462596
rect 247862 462476 247868 462528
rect 247920 462516 247926 462528
rect 427078 462516 427084 462528
rect 247920 462488 427084 462516
rect 247920 462476 247926 462488
rect 427078 462476 427084 462488
rect 427136 462476 427142 462528
rect 242802 462408 242808 462460
rect 242860 462448 242866 462460
rect 424318 462448 424324 462460
rect 242860 462420 424324 462448
rect 242860 462408 242866 462420
rect 424318 462408 424324 462420
rect 424376 462408 424382 462460
rect 3510 462340 3516 462392
rect 3568 462380 3574 462392
rect 370774 462380 370780 462392
rect 3568 462352 370780 462380
rect 3568 462340 3574 462352
rect 370774 462340 370780 462352
rect 370832 462340 370838 462392
rect 307294 461592 307300 461644
rect 307352 461632 307358 461644
rect 413278 461632 413284 461644
rect 307352 461604 413284 461632
rect 307352 461592 307358 461604
rect 413278 461592 413284 461604
rect 413336 461592 413342 461644
rect 236730 461388 236736 461440
rect 236788 461428 236794 461440
rect 373994 461428 374000 461440
rect 236788 461400 374000 461428
rect 236788 461388 236794 461400
rect 373994 461388 374000 461400
rect 374052 461388 374058 461440
rect 229738 461320 229744 461372
rect 229796 461360 229802 461372
rect 396074 461360 396080 461372
rect 229796 461332 396080 461360
rect 229796 461320 229802 461332
rect 396074 461320 396080 461332
rect 396132 461320 396138 461372
rect 250898 461252 250904 461304
rect 250956 461292 250962 461304
rect 417418 461292 417424 461304
rect 250956 461264 417424 461292
rect 250956 461252 250962 461264
rect 417418 461252 417424 461264
rect 417476 461252 417482 461304
rect 257246 461184 257252 461236
rect 257304 461224 257310 461236
rect 428458 461224 428464 461236
rect 257304 461196 428464 461224
rect 257304 461184 257310 461196
rect 428458 461184 428464 461196
rect 428516 461184 428522 461236
rect 228358 461116 228364 461168
rect 228416 461156 228422 461168
rect 400490 461156 400496 461168
rect 228416 461128 400496 461156
rect 228416 461116 228422 461128
rect 400490 461116 400496 461128
rect 400548 461116 400554 461168
rect 224218 461048 224224 461100
rect 224276 461088 224282 461100
rect 409874 461088 409880 461100
rect 224276 461060 409880 461088
rect 224276 461048 224282 461060
rect 409874 461048 409880 461060
rect 409932 461048 409938 461100
rect 269758 460980 269764 461032
rect 269816 461020 269822 461032
rect 567930 461020 567936 461032
rect 269816 460992 567936 461020
rect 269816 460980 269822 460992
rect 567930 460980 567936 460992
rect 567988 460980 567994 461032
rect 18690 460912 18696 460964
rect 18748 460952 18754 460964
rect 391106 460952 391112 460964
rect 18748 460924 391112 460952
rect 18748 460912 18754 460924
rect 391106 460912 391112 460924
rect 391164 460912 391170 460964
rect 201494 460844 201500 460896
rect 201552 460884 201558 460896
rect 331674 460884 331680 460896
rect 201552 460856 331680 460884
rect 201552 460844 201558 460856
rect 331674 460844 331680 460856
rect 331732 460844 331738 460896
rect 313182 460776 313188 460828
rect 313240 460816 313246 460828
rect 462314 460816 462320 460828
rect 313240 460788 462320 460816
rect 313240 460776 313246 460788
rect 462314 460776 462320 460788
rect 462372 460776 462378 460828
rect 315114 460708 315120 460760
rect 315172 460748 315178 460760
rect 477494 460748 477500 460760
rect 315172 460720 477500 460748
rect 315172 460708 315178 460720
rect 477494 460708 477500 460720
rect 477552 460708 477558 460760
rect 136634 460640 136640 460692
rect 136692 460680 136698 460692
rect 336366 460680 336372 460692
rect 136692 460652 336372 460680
rect 136692 460640 136698 460652
rect 336366 460640 336372 460652
rect 336424 460640 336430 460692
rect 308858 460572 308864 460624
rect 308916 460612 308922 460624
rect 527174 460612 527180 460624
rect 308916 460584 527180 460612
rect 308916 460572 308922 460584
rect 527174 460572 527180 460584
rect 527232 460572 527238 460624
rect 310422 460504 310428 460556
rect 310480 460544 310486 460556
rect 542354 460544 542360 460556
rect 310480 460516 542360 460544
rect 310480 460504 310486 460516
rect 542354 460504 542360 460516
rect 542412 460504 542418 460556
rect 71774 460436 71780 460488
rect 71832 460476 71838 460488
rect 341058 460476 341064 460488
rect 71832 460448 341064 460476
rect 71832 460436 71838 460448
rect 341058 460436 341064 460448
rect 341116 460436 341122 460488
rect 3602 460368 3608 460420
rect 3660 460408 3666 460420
rect 353570 460408 353576 460420
rect 3660 460380 353576 460408
rect 3660 460368 3666 460380
rect 353570 460368 353576 460380
rect 353628 460368 353634 460420
rect 3694 460300 3700 460352
rect 3752 460340 3758 460352
rect 358262 460340 358268 460352
rect 3752 460312 358268 460340
rect 3752 460300 3758 460312
rect 358262 460300 358268 460312
rect 358320 460300 358326 460352
rect 3786 460232 3792 460284
rect 3844 460272 3850 460284
rect 362954 460272 362960 460284
rect 3844 460244 362960 460272
rect 3844 460232 3850 460244
rect 362954 460232 362960 460244
rect 363012 460232 363018 460284
rect 3878 460164 3884 460216
rect 3936 460204 3942 460216
rect 367646 460204 367652 460216
rect 3936 460176 367652 460204
rect 3936 460164 3942 460176
rect 367646 460164 367652 460176
rect 367704 460164 367710 460216
rect 318242 460096 318248 460148
rect 318300 460136 318306 460148
rect 397454 460136 397460 460148
rect 318300 460108 397460 460136
rect 318300 460096 318306 460108
rect 397454 460096 397460 460108
rect 397512 460096 397518 460148
rect 266354 460028 266360 460080
rect 266412 460068 266418 460080
rect 327074 460068 327080 460080
rect 266412 460040 327080 460068
rect 266412 460028 266418 460040
rect 327074 460028 327080 460040
rect 327132 460028 327138 460080
rect 322842 459960 322848 460012
rect 322900 460000 322906 460012
rect 331214 460000 331220 460012
rect 322900 459972 331220 460000
rect 322900 459960 322906 459972
rect 331214 459960 331220 459972
rect 331272 459960 331278 460012
rect 282270 459552 282276 459604
rect 282328 459592 282334 459604
rect 308490 459592 308496 459604
rect 282328 459564 308496 459592
rect 282328 459552 282334 459564
rect 308490 459552 308496 459564
rect 308548 459552 308554 459604
rect 353294 459552 353300 459604
rect 353352 459592 353358 459604
rect 369210 459592 369216 459604
rect 353352 459564 369216 459592
rect 353352 459552 353358 459564
rect 369210 459552 369216 459564
rect 369268 459552 369274 459604
rect 235258 458872 235264 458924
rect 235316 458912 235322 458924
rect 377030 458912 377036 458924
rect 235316 458884 377036 458912
rect 235316 458872 235322 458884
rect 377030 458872 377036 458884
rect 377088 458872 377094 458924
rect 308490 458804 308496 458856
rect 308548 458844 308554 458856
rect 580350 458844 580356 458856
rect 308548 458816 580356 458844
rect 308548 458804 308554 458816
rect 580350 458804 580356 458816
rect 580408 458804 580414 458856
rect 274450 458736 274456 458788
rect 274508 458776 274514 458788
rect 416038 458776 416044 458788
rect 274508 458748 416044 458776
rect 274508 458736 274514 458748
rect 416038 458736 416044 458748
rect 416096 458736 416102 458788
rect 233970 458668 233976 458720
rect 234028 458708 234034 458720
rect 381722 458708 381728 458720
rect 234028 458680 381728 458708
rect 234028 458668 234034 458680
rect 381722 458668 381728 458680
rect 381780 458668 381786 458720
rect 232498 458600 232504 458652
rect 232556 458640 232562 458652
rect 386414 458640 386420 458652
rect 232556 458612 386420 458640
rect 232556 458600 232562 458612
rect 386414 458600 386420 458612
rect 386472 458600 386478 458652
rect 255682 458532 255688 458584
rect 255740 458572 255746 458584
rect 418798 458572 418804 458584
rect 255740 458544 418804 458572
rect 255740 458532 255746 458544
rect 418798 458532 418804 458544
rect 418856 458532 418862 458584
rect 266262 458464 266268 458516
rect 266320 458504 266326 458516
rect 431218 458504 431224 458516
rect 266320 458476 431224 458504
rect 266320 458464 266326 458476
rect 431218 458464 431224 458476
rect 431276 458464 431282 458516
rect 246298 458396 246304 458448
rect 246356 458436 246362 458448
rect 414658 458436 414664 458448
rect 246356 458408 414664 458436
rect 246356 458396 246362 458408
rect 414658 458396 414664 458408
rect 414716 458396 414722 458448
rect 225598 458328 225604 458380
rect 225656 458368 225662 458380
rect 405182 458368 405188 458380
rect 225656 458340 405188 458368
rect 225656 458328 225662 458340
rect 405182 458328 405188 458340
rect 405240 458328 405246 458380
rect 241422 458260 241428 458312
rect 241480 458300 241486 458312
rect 580258 458300 580264 458312
rect 241480 458272 580264 458300
rect 241480 458260 241486 458272
rect 580258 458260 580264 458272
rect 580316 458260 580322 458312
rect 3418 458192 3424 458244
rect 3476 458232 3482 458244
rect 372660 458232 372666 458244
rect 3476 458204 372666 458232
rect 3476 458192 3482 458204
rect 372660 458192 372666 458204
rect 372718 458192 372724 458244
rect 273226 457592 292574 457620
rect 238018 457512 238024 457564
rect 238076 457552 238082 457564
rect 239398 457552 239404 457564
rect 238076 457524 239404 457552
rect 238076 457512 238082 457524
rect 239398 457512 239404 457524
rect 239456 457512 239462 457564
rect 3510 457444 3516 457496
rect 3568 457484 3574 457496
rect 273226 457484 273254 457592
rect 280126 457524 289814 457552
rect 3568 457456 273254 457484
rect 3568 457444 3574 457456
rect 275922 457444 275928 457496
rect 275980 457484 275986 457496
rect 280126 457484 280154 457524
rect 275980 457456 280154 457484
rect 275980 457444 275986 457456
rect 283650 457444 283656 457496
rect 283708 457444 283714 457496
rect 283668 456804 283696 457444
rect 289786 457280 289814 457524
rect 292546 457484 292574 457592
rect 353294 457484 353300 457496
rect 292546 457456 353300 457484
rect 353294 457444 353300 457456
rect 353352 457444 353358 457496
rect 412082 457444 412088 457496
rect 412140 457484 412146 457496
rect 414106 457484 414112 457496
rect 412140 457456 414112 457484
rect 412140 457444 412146 457456
rect 414106 457444 414112 457456
rect 414164 457444 414170 457496
rect 289786 457252 292574 457280
rect 292546 456872 292574 457252
rect 432598 456872 432604 456884
rect 292546 456844 432604 456872
rect 432598 456832 432604 456844
rect 432656 456832 432662 456884
rect 580166 456804 580172 456816
rect 283668 456776 580172 456804
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 457438 431876 457444 431928
rect 457496 431916 457502 431928
rect 579614 431916 579620 431928
rect 457496 431888 579620 431916
rect 457496 431876 457502 431888
rect 579614 431876 579620 431888
rect 579672 431876 579678 431928
rect 3418 411204 3424 411256
rect 3476 411244 3482 411256
rect 235350 411244 235356 411256
rect 3476 411216 235356 411244
rect 3476 411204 3482 411216
rect 235350 411204 235356 411216
rect 235408 411204 235414 411256
rect 454678 405628 454684 405680
rect 454736 405668 454742 405680
rect 579614 405668 579620 405680
rect 454736 405640 579620 405668
rect 454736 405628 454742 405640
rect 579614 405628 579620 405640
rect 579672 405628 579678 405680
rect 3234 398760 3240 398812
rect 3292 398800 3298 398812
rect 235902 398800 235908 398812
rect 3292 398772 235908 398800
rect 3292 398760 3298 398772
rect 235902 398760 235908 398772
rect 235960 398760 235966 398812
rect 432598 379448 432604 379500
rect 432656 379488 432662 379500
rect 580166 379488 580172 379500
rect 432656 379460 580172 379488
rect 432656 379448 432662 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 3234 372512 3240 372564
rect 3292 372552 3298 372564
rect 235258 372552 235264 372564
rect 3292 372524 235264 372552
rect 3292 372512 3298 372524
rect 235258 372512 235264 372524
rect 235316 372512 235322 372564
rect 435358 365644 435364 365696
rect 435416 365684 435422 365696
rect 580166 365684 580172 365696
rect 435416 365656 580172 365684
rect 435416 365644 435422 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 3326 358708 3332 358760
rect 3384 358748 3390 358760
rect 215938 358748 215944 358760
rect 3384 358720 215944 358748
rect 3384 358708 3390 358720
rect 215938 358708 215944 358720
rect 215996 358708 216002 358760
rect 416038 353200 416044 353252
rect 416096 353240 416102 353252
rect 580166 353240 580172 353252
rect 416096 353212 580172 353240
rect 416096 353200 416102 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 3142 346332 3148 346384
rect 3200 346372 3206 346384
rect 13078 346372 13084 346384
rect 3200 346344 13084 346372
rect 3200 346332 3206 346344
rect 13078 346332 13084 346344
rect 13136 346332 13142 346384
rect 256050 336676 256056 336728
rect 256108 336716 256114 336728
rect 257798 336716 257804 336728
rect 256108 336688 257804 336716
rect 256108 336676 256114 336688
rect 257798 336676 257804 336688
rect 257856 336676 257862 336728
rect 264238 336676 264244 336728
rect 264296 336716 264302 336728
rect 266354 336716 266360 336728
rect 264296 336688 266360 336716
rect 264296 336676 264302 336688
rect 266354 336676 266360 336688
rect 266412 336676 266418 336728
rect 271138 336676 271144 336728
rect 271196 336716 271202 336728
rect 273254 336716 273260 336728
rect 271196 336688 273260 336716
rect 271196 336676 271202 336688
rect 273254 336676 273260 336688
rect 273312 336676 273318 336728
rect 273898 336676 273904 336728
rect 273956 336716 273962 336728
rect 275002 336716 275008 336728
rect 273956 336688 275008 336716
rect 273956 336676 273962 336688
rect 275002 336676 275008 336688
rect 275060 336676 275066 336728
rect 278866 336676 278872 336728
rect 278924 336716 278930 336728
rect 279142 336716 279148 336728
rect 278924 336688 279148 336716
rect 278924 336676 278930 336688
rect 279142 336676 279148 336688
rect 279200 336676 279206 336728
rect 279418 336676 279424 336728
rect 279476 336716 279482 336728
rect 280430 336716 280436 336728
rect 279476 336688 280436 336716
rect 279476 336676 279482 336688
rect 280430 336676 280436 336688
rect 280488 336676 280494 336728
rect 284478 336676 284484 336728
rect 284536 336716 284542 336728
rect 284846 336716 284852 336728
rect 284536 336688 284852 336716
rect 284536 336676 284542 336688
rect 284846 336676 284852 336688
rect 284904 336676 284910 336728
rect 287698 336676 287704 336728
rect 287756 336716 287762 336728
rect 288986 336716 288992 336728
rect 287756 336688 288992 336716
rect 287756 336676 287762 336688
rect 288986 336676 288992 336688
rect 289044 336676 289050 336728
rect 289170 336676 289176 336728
rect 289228 336716 289234 336728
rect 290366 336716 290372 336728
rect 289228 336688 290372 336716
rect 289228 336676 289234 336688
rect 290366 336676 290372 336688
rect 290424 336676 290430 336728
rect 293218 336676 293224 336728
rect 293276 336716 293282 336728
rect 294230 336716 294236 336728
rect 293276 336688 294236 336716
rect 293276 336676 293282 336688
rect 294230 336676 294236 336688
rect 294288 336676 294294 336728
rect 296806 336676 296812 336728
rect 296864 336716 296870 336728
rect 297542 336716 297548 336728
rect 296864 336688 297548 336716
rect 296864 336676 296870 336688
rect 297542 336676 297548 336688
rect 297600 336676 297606 336728
rect 298738 336676 298744 336728
rect 298796 336716 298802 336728
rect 300026 336716 300032 336728
rect 298796 336688 300032 336716
rect 298796 336676 298802 336688
rect 300026 336676 300032 336688
rect 300084 336676 300090 336728
rect 300854 336676 300860 336728
rect 300912 336716 300918 336728
rect 301130 336716 301136 336728
rect 300912 336688 301136 336716
rect 300912 336676 300918 336688
rect 301130 336676 301136 336688
rect 301188 336676 301194 336728
rect 302234 336676 302240 336728
rect 302292 336716 302298 336728
rect 302510 336716 302516 336728
rect 302292 336688 302516 336716
rect 302292 336676 302298 336688
rect 302510 336676 302516 336688
rect 302568 336676 302574 336728
rect 303614 336676 303620 336728
rect 303672 336716 303678 336728
rect 303982 336716 303988 336728
rect 303672 336688 303988 336716
rect 303672 336676 303678 336688
rect 303982 336676 303988 336688
rect 304040 336676 304046 336728
rect 309870 336676 309876 336728
rect 309928 336716 309934 336728
rect 312722 336716 312728 336728
rect 309928 336688 312728 336716
rect 309928 336676 309934 336688
rect 312722 336676 312728 336688
rect 312780 336676 312786 336728
rect 318886 336676 318892 336728
rect 318944 336716 318950 336728
rect 319070 336716 319076 336728
rect 318944 336688 319076 336716
rect 318944 336676 318950 336688
rect 319070 336676 319076 336688
rect 319128 336676 319134 336728
rect 327718 336676 327724 336728
rect 327776 336716 327782 336728
rect 331214 336716 331220 336728
rect 327776 336688 331220 336716
rect 327776 336676 327782 336688
rect 331214 336676 331220 336688
rect 331272 336676 331278 336728
rect 334066 336676 334072 336728
rect 334124 336716 334130 336728
rect 334342 336716 334348 336728
rect 334124 336688 334348 336716
rect 334124 336676 334130 336688
rect 334342 336676 334348 336688
rect 334400 336676 334406 336728
rect 336734 336676 336740 336728
rect 336792 336716 336798 336728
rect 337102 336716 337108 336728
rect 336792 336688 337108 336716
rect 336792 336676 336798 336688
rect 337102 336676 337108 336688
rect 337160 336676 337166 336728
rect 348602 336676 348608 336728
rect 348660 336716 348666 336728
rect 349798 336716 349804 336728
rect 348660 336688 349804 336716
rect 348660 336676 348666 336688
rect 349798 336676 349804 336688
rect 349856 336676 349862 336728
rect 353478 336676 353484 336728
rect 353536 336716 353542 336728
rect 353662 336716 353668 336728
rect 353536 336688 353668 336716
rect 353536 336676 353542 336688
rect 353662 336676 353668 336688
rect 353720 336676 353726 336728
rect 356238 336676 356244 336728
rect 356296 336716 356302 336728
rect 356422 336716 356428 336728
rect 356296 336688 356428 336716
rect 356296 336676 356302 336688
rect 356422 336676 356428 336688
rect 356480 336676 356486 336728
rect 372706 336676 372712 336728
rect 372764 336716 372770 336728
rect 372982 336716 372988 336728
rect 372764 336688 372988 336716
rect 372764 336676 372770 336688
rect 372982 336676 372988 336688
rect 373040 336676 373046 336728
rect 376202 336676 376208 336728
rect 376260 336716 376266 336728
rect 377398 336716 377404 336728
rect 376260 336688 377404 336716
rect 376260 336676 376266 336688
rect 377398 336676 377404 336688
rect 377456 336676 377462 336728
rect 378318 336676 378324 336728
rect 378376 336716 378382 336728
rect 378502 336716 378508 336728
rect 378376 336688 378508 336716
rect 378376 336676 378382 336688
rect 378502 336676 378508 336688
rect 378560 336676 378566 336728
rect 386598 336676 386604 336728
rect 386656 336716 386662 336728
rect 386782 336716 386788 336728
rect 386656 336688 386788 336716
rect 386656 336676 386662 336688
rect 386782 336676 386788 336688
rect 386840 336676 386846 336728
rect 256142 336608 256148 336660
rect 256200 336648 256206 336660
rect 260834 336648 260840 336660
rect 256200 336620 260840 336648
rect 256200 336608 256206 336620
rect 260834 336608 260840 336620
rect 260892 336608 260898 336660
rect 268378 336608 268384 336660
rect 268436 336648 268442 336660
rect 272150 336648 272156 336660
rect 268436 336620 272156 336648
rect 268436 336608 268442 336620
rect 272150 336608 272156 336620
rect 272208 336608 272214 336660
rect 303522 336608 303528 336660
rect 303580 336648 303586 336660
rect 311894 336648 311900 336660
rect 303580 336620 311900 336648
rect 303580 336608 303586 336620
rect 311894 336608 311900 336620
rect 311952 336608 311958 336660
rect 318058 336608 318064 336660
rect 318116 336648 318122 336660
rect 320450 336648 320456 336660
rect 318116 336620 320456 336648
rect 318116 336608 318122 336620
rect 320450 336608 320456 336620
rect 320508 336608 320514 336660
rect 257338 336540 257344 336592
rect 257396 336580 257402 336592
rect 268838 336580 268844 336592
rect 257396 336552 268844 336580
rect 257396 336540 257402 336552
rect 268838 336540 268844 336552
rect 268896 336540 268902 336592
rect 305730 336540 305736 336592
rect 305788 336580 305794 336592
rect 316034 336580 316040 336592
rect 305788 336552 316040 336580
rect 305788 336540 305794 336552
rect 316034 336540 316040 336552
rect 316092 336540 316098 336592
rect 316678 336540 316684 336592
rect 316736 336580 316742 336592
rect 322106 336580 322112 336592
rect 316736 336552 322112 336580
rect 316736 336540 316742 336552
rect 322106 336540 322112 336552
rect 322164 336540 322170 336592
rect 348694 336540 348700 336592
rect 348752 336580 348758 336592
rect 370498 336580 370504 336592
rect 348752 336552 370504 336580
rect 348752 336540 348758 336552
rect 370498 336540 370504 336552
rect 370556 336540 370562 336592
rect 377490 336540 377496 336592
rect 377548 336580 377554 336592
rect 399478 336580 399484 336592
rect 377548 336552 399484 336580
rect 377548 336540 377554 336552
rect 399478 336540 399484 336552
rect 399536 336540 399542 336592
rect 233878 336472 233884 336524
rect 233936 336512 233942 336524
rect 264698 336512 264704 336524
rect 233936 336484 264704 336512
rect 233936 336472 233942 336484
rect 264698 336472 264704 336484
rect 264756 336472 264762 336524
rect 307018 336472 307024 336524
rect 307076 336512 307082 336524
rect 322934 336512 322940 336524
rect 307076 336484 322940 336512
rect 307076 336472 307082 336484
rect 322934 336472 322940 336484
rect 322992 336472 322998 336524
rect 323578 336472 323584 336524
rect 323636 336512 323642 336524
rect 324590 336512 324596 336524
rect 323636 336484 324596 336512
rect 323636 336472 323642 336484
rect 324590 336472 324596 336484
rect 324648 336472 324654 336524
rect 344278 336472 344284 336524
rect 344336 336512 344342 336524
rect 359550 336512 359556 336524
rect 344336 336484 359556 336512
rect 344336 336472 344342 336484
rect 359550 336472 359556 336484
rect 359608 336472 359614 336524
rect 370774 336472 370780 336524
rect 370832 336512 370838 336524
rect 395338 336512 395344 336524
rect 370832 336484 395344 336512
rect 370832 336472 370838 336484
rect 395338 336472 395344 336484
rect 395396 336472 395402 336524
rect 255958 336404 255964 336456
rect 256016 336444 256022 336456
rect 296162 336444 296168 336456
rect 256016 336416 296168 336444
rect 256016 336404 256022 336416
rect 296162 336404 296168 336416
rect 296220 336404 296226 336456
rect 301498 336404 301504 336456
rect 301556 336444 301562 336456
rect 317690 336444 317696 336456
rect 301556 336416 317696 336444
rect 301556 336404 301562 336416
rect 317690 336404 317696 336416
rect 317748 336404 317754 336456
rect 342070 336404 342076 336456
rect 342128 336444 342134 336456
rect 363598 336444 363604 336456
rect 342128 336416 363604 336444
rect 342128 336404 342134 336416
rect 363598 336404 363604 336416
rect 363656 336404 363662 336456
rect 369946 336404 369952 336456
rect 370004 336444 370010 336456
rect 396718 336444 396724 336456
rect 370004 336416 396724 336444
rect 370004 336404 370010 336416
rect 396718 336404 396724 336416
rect 396776 336404 396782 336456
rect 243538 336336 243544 336388
rect 243596 336376 243602 336388
rect 287882 336376 287888 336388
rect 243596 336348 287888 336376
rect 243596 336336 243602 336348
rect 287882 336336 287888 336348
rect 287940 336336 287946 336388
rect 305638 336336 305644 336388
rect 305696 336376 305702 336388
rect 323486 336376 323492 336388
rect 305696 336348 323492 336376
rect 305696 336336 305702 336348
rect 323486 336336 323492 336348
rect 323544 336336 323550 336388
rect 346762 336336 346768 336388
rect 346820 336376 346826 336388
rect 378778 336376 378784 336388
rect 346820 336348 378784 336376
rect 346820 336336 346826 336348
rect 378778 336336 378784 336348
rect 378836 336336 378842 336388
rect 382366 336336 382372 336388
rect 382424 336376 382430 336388
rect 407758 336376 407764 336388
rect 382424 336348 407764 336376
rect 382424 336336 382430 336348
rect 407758 336336 407764 336348
rect 407816 336336 407822 336388
rect 242158 336268 242164 336320
rect 242216 336308 242222 336320
rect 296438 336308 296444 336320
rect 242216 336280 296444 336308
rect 242216 336268 242222 336280
rect 296438 336268 296444 336280
rect 296496 336268 296502 336320
rect 304258 336268 304264 336320
rect 304316 336308 304322 336320
rect 322658 336308 322664 336320
rect 304316 336280 322664 336308
rect 304316 336268 304322 336280
rect 322658 336268 322664 336280
rect 322716 336268 322722 336320
rect 340046 336268 340052 336320
rect 340104 336308 340110 336320
rect 341518 336308 341524 336320
rect 340104 336280 341524 336308
rect 340104 336268 340110 336280
rect 341518 336268 341524 336280
rect 341576 336268 341582 336320
rect 345106 336268 345112 336320
rect 345164 336308 345170 336320
rect 371878 336308 371884 336320
rect 345164 336280 371884 336308
rect 345164 336268 345170 336280
rect 371878 336268 371884 336280
rect 371936 336268 371942 336320
rect 374270 336268 374276 336320
rect 374328 336308 374334 336320
rect 410518 336308 410524 336320
rect 374328 336280 410524 336308
rect 374328 336268 374334 336280
rect 410518 336268 410524 336280
rect 410576 336268 410582 336320
rect 247678 336200 247684 336252
rect 247736 336240 247742 336252
rect 307754 336240 307760 336252
rect 247736 336212 307760 336240
rect 247736 336200 247742 336212
rect 307754 336200 307760 336212
rect 307812 336200 307818 336252
rect 309778 336200 309784 336252
rect 309836 336240 309842 336252
rect 320174 336240 320180 336252
rect 309836 336212 320180 336240
rect 309836 336200 309842 336212
rect 320174 336200 320180 336212
rect 320232 336200 320238 336252
rect 322198 336200 322204 336252
rect 322256 336240 322262 336252
rect 330938 336240 330944 336252
rect 322256 336212 330944 336240
rect 322256 336200 322262 336212
rect 330938 336200 330944 336212
rect 330996 336200 331002 336252
rect 340138 336200 340144 336252
rect 340196 336240 340202 336252
rect 356054 336240 356060 336252
rect 340196 336212 356060 336240
rect 340196 336200 340202 336212
rect 356054 336200 356060 336212
rect 356112 336200 356118 336252
rect 358906 336200 358912 336252
rect 358964 336240 358970 336252
rect 436094 336240 436100 336252
rect 358964 336212 436100 336240
rect 358964 336200 358970 336212
rect 436094 336200 436100 336212
rect 436152 336200 436158 336252
rect 117314 336132 117320 336184
rect 117372 336172 117378 336184
rect 284294 336172 284300 336184
rect 117372 336144 284300 336172
rect 117372 336132 117378 336144
rect 284294 336132 284300 336144
rect 284352 336132 284358 336184
rect 297542 336132 297548 336184
rect 297600 336172 297606 336184
rect 298646 336172 298652 336184
rect 297600 336144 298652 336172
rect 297600 336132 297606 336144
rect 298646 336132 298652 336144
rect 298704 336132 298710 336184
rect 300118 336132 300124 336184
rect 300176 336172 300182 336184
rect 321830 336172 321836 336184
rect 300176 336144 321836 336172
rect 300176 336132 300182 336144
rect 321830 336132 321836 336144
rect 321888 336132 321894 336184
rect 360562 336132 360568 336184
rect 360620 336172 360626 336184
rect 442994 336172 443000 336184
rect 360620 336144 443000 336172
rect 360620 336132 360626 336144
rect 442994 336132 443000 336144
rect 443052 336132 443058 336184
rect 110414 336064 110420 336116
rect 110472 336104 110478 336116
rect 282638 336104 282644 336116
rect 110472 336076 282644 336104
rect 110472 336064 110478 336076
rect 282638 336064 282644 336076
rect 282696 336064 282702 336116
rect 295978 336064 295984 336116
rect 296036 336104 296042 336116
rect 319346 336104 319352 336116
rect 296036 336076 319352 336104
rect 296036 336064 296042 336076
rect 319346 336064 319352 336076
rect 319404 336064 319410 336116
rect 320818 336064 320824 336116
rect 320876 336104 320882 336116
rect 330110 336104 330116 336116
rect 320876 336076 330116 336104
rect 320876 336064 320882 336076
rect 330110 336064 330116 336076
rect 330168 336064 330174 336116
rect 342346 336064 342352 336116
rect 342404 336104 342410 336116
rect 360838 336104 360844 336116
rect 342404 336076 360844 336104
rect 342404 336064 342410 336076
rect 360838 336064 360844 336076
rect 360896 336064 360902 336116
rect 362218 336064 362224 336116
rect 362276 336104 362282 336116
rect 449894 336104 449900 336116
rect 362276 336076 449900 336104
rect 362276 336064 362282 336076
rect 449894 336064 449900 336076
rect 449952 336064 449958 336116
rect 10318 335996 10324 336048
rect 10376 336036 10382 336048
rect 10376 336008 238754 336036
rect 10376 335996 10382 336008
rect 238726 335968 238754 336008
rect 269758 335996 269764 336048
rect 269816 336036 269822 336048
rect 271046 336036 271052 336048
rect 269816 336008 271052 336036
rect 269816 335996 269822 336008
rect 271046 335996 271052 336008
rect 271104 335996 271110 336048
rect 285674 335996 285680 336048
rect 285732 336036 285738 336048
rect 294506 336036 294512 336048
rect 285732 336008 294512 336036
rect 285732 335996 285738 336008
rect 294506 335996 294512 336008
rect 294564 335996 294570 336048
rect 297174 335996 297180 336048
rect 297232 336036 297238 336048
rect 324314 336036 324320 336048
rect 297232 336008 324320 336036
rect 297232 335996 297238 336008
rect 324314 335996 324320 336008
rect 324372 335996 324378 336048
rect 341242 335996 341248 336048
rect 341300 336036 341306 336048
rect 359458 336036 359464 336048
rect 341300 336008 359464 336036
rect 341300 335996 341306 336008
rect 359458 335996 359464 336008
rect 359516 335996 359522 336048
rect 363874 335996 363880 336048
rect 363932 336036 363938 336048
rect 456794 336036 456800 336048
rect 363932 336008 456800 336036
rect 363932 335996 363938 336008
rect 456794 335996 456800 336008
rect 456852 335996 456858 336048
rect 258350 335968 258356 335980
rect 238726 335940 258356 335968
rect 258350 335928 258356 335940
rect 258408 335928 258414 335980
rect 284294 335928 284300 335980
rect 284352 335968 284358 335980
rect 286226 335968 286232 335980
rect 284352 335940 286232 335968
rect 284352 335928 284358 335940
rect 286226 335928 286232 335940
rect 286284 335928 286290 335980
rect 293310 335928 293316 335980
rect 293368 335968 293374 335980
rect 293954 335968 293960 335980
rect 293368 335940 293960 335968
rect 293368 335928 293374 335940
rect 293954 335928 293960 335940
rect 294012 335928 294018 335980
rect 356698 335860 356704 335912
rect 356756 335900 356762 335912
rect 360562 335900 360568 335912
rect 356756 335872 360568 335900
rect 356756 335860 356762 335872
rect 360562 335860 360568 335872
rect 360620 335860 360626 335912
rect 365806 335860 365812 335912
rect 365864 335900 365870 335912
rect 369118 335900 369124 335912
rect 365864 335872 369124 335900
rect 365864 335860 365870 335872
rect 369118 335860 369124 335872
rect 369176 335860 369182 335912
rect 271230 335792 271236 335844
rect 271288 335832 271294 335844
rect 272978 335832 272984 335844
rect 271288 335804 272984 335832
rect 271288 335792 271294 335804
rect 272978 335792 272984 335804
rect 273036 335792 273042 335844
rect 343726 335792 343732 335844
rect 343784 335832 343790 335844
rect 345658 335832 345664 335844
rect 343784 335804 345664 335832
rect 343784 335792 343790 335804
rect 345658 335792 345664 335804
rect 345716 335792 345722 335844
rect 357526 335724 357532 335776
rect 357584 335764 357590 335776
rect 360930 335764 360936 335776
rect 357584 335736 360936 335764
rect 357584 335724 357590 335736
rect 360930 335724 360936 335736
rect 360988 335724 360994 335776
rect 261478 335656 261484 335708
rect 261536 335696 261542 335708
rect 263042 335696 263048 335708
rect 261536 335668 263048 335696
rect 261536 335656 261542 335668
rect 263042 335656 263048 335668
rect 263100 335656 263106 335708
rect 275278 335656 275284 335708
rect 275336 335696 275342 335708
rect 276290 335696 276296 335708
rect 275336 335668 276296 335696
rect 275336 335656 275342 335668
rect 276290 335656 276296 335668
rect 276348 335656 276354 335708
rect 287790 335656 287796 335708
rect 287848 335696 287854 335708
rect 288710 335696 288716 335708
rect 287848 335668 288716 335696
rect 287848 335656 287854 335668
rect 288710 335656 288716 335668
rect 288768 335656 288774 335708
rect 291838 335656 291844 335708
rect 291896 335696 291902 335708
rect 293126 335696 293132 335708
rect 291896 335668 293132 335696
rect 291896 335656 291902 335668
rect 293126 335656 293132 335668
rect 293184 335656 293190 335708
rect 315298 335656 315304 335708
rect 315356 335696 315362 335708
rect 317138 335696 317144 335708
rect 315356 335668 317144 335696
rect 315356 335656 315362 335668
rect 317138 335656 317144 335668
rect 317196 335656 317202 335708
rect 361666 335656 361672 335708
rect 361724 335696 361730 335708
rect 363690 335696 363696 335708
rect 361724 335668 363696 335696
rect 361724 335656 361730 335668
rect 363690 335656 363696 335668
rect 363748 335656 363754 335708
rect 297450 335588 297456 335640
rect 297508 335628 297514 335640
rect 298094 335628 298100 335640
rect 297508 335600 298100 335628
rect 297508 335588 297514 335600
rect 298094 335588 298100 335600
rect 298152 335588 298158 335640
rect 289078 335520 289084 335572
rect 289136 335560 289142 335572
rect 289814 335560 289820 335572
rect 289136 335532 289820 335560
rect 289136 335520 289142 335532
rect 289814 335520 289820 335532
rect 289872 335520 289878 335572
rect 296162 335452 296168 335504
rect 296220 335492 296226 335504
rect 298370 335492 298376 335504
rect 296220 335464 298376 335492
rect 296220 335452 296226 335464
rect 298370 335452 298376 335464
rect 298428 335452 298434 335504
rect 311158 335452 311164 335504
rect 311216 335492 311222 335504
rect 317966 335492 317972 335504
rect 311216 335464 317972 335492
rect 311216 335452 311222 335464
rect 317966 335452 317972 335464
rect 318024 335452 318030 335504
rect 296070 335384 296076 335436
rect 296128 335424 296134 335436
rect 297266 335424 297272 335436
rect 296128 335396 297272 335424
rect 296128 335384 296134 335396
rect 297266 335384 297272 335396
rect 297324 335384 297330 335436
rect 323670 335384 323676 335436
rect 323728 335424 323734 335436
rect 326798 335424 326804 335436
rect 323728 335396 326804 335424
rect 323728 335384 323734 335396
rect 326798 335384 326804 335396
rect 326856 335384 326862 335436
rect 392026 335384 392032 335436
rect 392084 335424 392090 335436
rect 393958 335424 393964 335436
rect 392084 335396 393964 335424
rect 392084 335384 392090 335396
rect 393958 335384 393964 335396
rect 394016 335384 394022 335436
rect 257430 335316 257436 335368
rect 257488 335356 257494 335368
rect 259178 335356 259184 335368
rect 257488 335328 259184 335356
rect 257488 335316 257494 335328
rect 259178 335316 259184 335328
rect 259236 335316 259242 335368
rect 286318 335316 286324 335368
rect 286376 335356 286382 335368
rect 287606 335356 287612 335368
rect 286376 335328 287612 335356
rect 286376 335316 286382 335328
rect 287606 335316 287612 335328
rect 287664 335316 287670 335368
rect 296254 335316 296260 335368
rect 296312 335356 296318 335368
rect 296990 335356 296996 335368
rect 296312 335328 296996 335356
rect 296312 335316 296318 335328
rect 296990 335316 296996 335328
rect 297048 335316 297054 335368
rect 302878 335316 302884 335368
rect 302936 335356 302942 335368
rect 306650 335356 306656 335368
rect 302936 335328 306656 335356
rect 302936 335316 302942 335328
rect 306650 335316 306656 335328
rect 306708 335316 306714 335368
rect 313918 335316 313924 335368
rect 313976 335356 313982 335368
rect 316862 335356 316868 335368
rect 313976 335328 316868 335356
rect 313976 335316 313982 335328
rect 316862 335316 316868 335328
rect 316920 335316 316926 335368
rect 324958 335316 324964 335368
rect 325016 335356 325022 335368
rect 325970 335356 325976 335368
rect 325016 335328 325976 335356
rect 325016 335316 325022 335328
rect 325970 335316 325976 335328
rect 326028 335316 326034 335368
rect 283190 335248 283196 335300
rect 283248 335288 283254 335300
rect 283374 335288 283380 335300
rect 283248 335260 283380 335288
rect 283248 335248 283254 335260
rect 283374 335248 283380 335260
rect 283432 335248 283438 335300
rect 332870 335248 332876 335300
rect 332928 335288 332934 335300
rect 333054 335288 333060 335300
rect 332928 335260 333060 335288
rect 332928 335248 332934 335260
rect 333054 335248 333060 335260
rect 333112 335248 333118 335300
rect 234614 334772 234620 334824
rect 234672 334812 234678 334824
rect 303522 334812 303528 334824
rect 234672 334784 303528 334812
rect 234672 334772 234678 334784
rect 303522 334772 303528 334784
rect 303580 334772 303586 334824
rect 205634 334704 205640 334756
rect 205692 334744 205698 334756
rect 304994 334744 305000 334756
rect 205692 334716 305000 334744
rect 205692 334704 205698 334716
rect 304994 334704 305000 334716
rect 305052 334704 305058 334756
rect 359366 334704 359372 334756
rect 359424 334744 359430 334756
rect 438854 334744 438860 334756
rect 359424 334716 438860 334744
rect 359424 334704 359430 334716
rect 438854 334704 438860 334716
rect 438912 334704 438918 334756
rect 160094 334636 160100 334688
rect 160152 334676 160158 334688
rect 285674 334676 285680 334688
rect 160152 334648 285680 334676
rect 160152 334636 160158 334648
rect 285674 334636 285680 334648
rect 285732 334636 285738 334688
rect 369210 334636 369216 334688
rect 369268 334676 369274 334688
rect 480254 334676 480260 334688
rect 369268 334648 480260 334676
rect 369268 334636 369274 334648
rect 480254 334636 480260 334648
rect 480312 334636 480318 334688
rect 14458 334568 14464 334620
rect 14516 334608 14522 334620
rect 259822 334608 259828 334620
rect 14516 334580 259828 334608
rect 14516 334568 14522 334580
rect 259822 334568 259828 334580
rect 259880 334568 259886 334620
rect 380802 334568 380808 334620
rect 380860 334608 380866 334620
rect 529934 334608 529940 334620
rect 380860 334580 529940 334608
rect 380860 334568 380866 334580
rect 529934 334568 529940 334580
rect 529992 334568 529998 334620
rect 248414 333412 248420 333464
rect 248472 333452 248478 333464
rect 314930 333452 314936 333464
rect 248472 333424 314936 333452
rect 248472 333412 248478 333424
rect 314930 333412 314936 333424
rect 314988 333412 314994 333464
rect 220814 333344 220820 333396
rect 220872 333384 220878 333396
rect 308582 333384 308588 333396
rect 220872 333356 308588 333384
rect 220872 333344 220878 333356
rect 308582 333344 308588 333356
rect 308640 333344 308646 333396
rect 360470 333344 360476 333396
rect 360528 333384 360534 333396
rect 441614 333384 441620 333396
rect 360528 333356 441620 333384
rect 360528 333344 360534 333356
rect 441614 333344 441620 333356
rect 441672 333344 441678 333396
rect 125594 333276 125600 333328
rect 125652 333316 125658 333328
rect 284294 333316 284300 333328
rect 125652 333288 284300 333316
rect 125652 333276 125658 333288
rect 284294 333276 284300 333288
rect 284352 333276 284358 333328
rect 494054 333316 494060 333328
rect 373966 333288 494060 333316
rect 13078 333208 13084 333260
rect 13136 333248 13142 333260
rect 13136 333220 238754 333248
rect 13136 333208 13142 333220
rect 238726 333180 238754 333220
rect 258626 333180 258632 333192
rect 238726 333152 258632 333180
rect 258626 333140 258632 333152
rect 258684 333140 258690 333192
rect 372522 333072 372528 333124
rect 372580 333112 372586 333124
rect 373966 333112 373994 333288
rect 494054 333276 494060 333288
rect 494112 333276 494118 333328
rect 384942 333208 384948 333260
rect 385000 333248 385006 333260
rect 547874 333248 547880 333260
rect 385000 333220 547880 333248
rect 385000 333208 385006 333220
rect 547874 333208 547880 333220
rect 547932 333208 547938 333260
rect 372580 333084 373994 333112
rect 372580 333072 372586 333084
rect 242894 331984 242900 332036
rect 242952 332024 242958 332036
rect 313826 332024 313832 332036
rect 242952 331996 313832 332024
rect 242952 331984 242958 331996
rect 313826 331984 313832 331996
rect 313884 331984 313890 332036
rect 349614 331984 349620 332036
rect 349672 332024 349678 332036
rect 396074 332024 396080 332036
rect 349672 331996 396080 332024
rect 349672 331984 349678 331996
rect 396074 331984 396080 331996
rect 396132 331984 396138 332036
rect 207014 331916 207020 331968
rect 207072 331956 207078 331968
rect 305362 331956 305368 331968
rect 207072 331928 305368 331956
rect 207072 331916 207078 331928
rect 305362 331916 305368 331928
rect 305420 331916 305426 331968
rect 371694 331916 371700 331968
rect 371752 331956 371758 331968
rect 489914 331956 489920 331968
rect 371752 331928 489920 331956
rect 371752 331916 371758 331928
rect 489914 331916 489920 331928
rect 489972 331916 489978 331968
rect 97994 331848 98000 331900
rect 98052 331888 98058 331900
rect 279878 331888 279884 331900
rect 98052 331860 279884 331888
rect 98052 331848 98058 331860
rect 279878 331848 279884 331860
rect 279936 331848 279942 331900
rect 384206 331848 384212 331900
rect 384264 331888 384270 331900
rect 543734 331888 543740 331900
rect 384264 331860 543740 331888
rect 384264 331848 384270 331860
rect 543734 331848 543740 331860
rect 543792 331848 543798 331900
rect 377030 331168 377036 331220
rect 377088 331208 377094 331220
rect 377214 331208 377220 331220
rect 377088 331180 377220 331208
rect 377088 331168 377094 331180
rect 377214 331168 377220 331180
rect 377272 331168 377278 331220
rect 327350 330896 327356 330948
rect 327408 330896 327414 330948
rect 292758 330692 292764 330744
rect 292816 330732 292822 330744
rect 292942 330732 292948 330744
rect 292816 330704 292948 330732
rect 292816 330692 292822 330704
rect 292942 330692 292948 330704
rect 293000 330692 293006 330744
rect 253934 330624 253940 330676
rect 253992 330664 253998 330676
rect 316310 330664 316316 330676
rect 253992 330636 316316 330664
rect 253992 330624 253998 330636
rect 316310 330624 316316 330636
rect 316368 330624 316374 330676
rect 327368 330608 327396 330896
rect 334342 330760 334348 330812
rect 334400 330760 334406 330812
rect 334360 330608 334388 330760
rect 352006 330624 352012 330676
rect 352064 330664 352070 330676
rect 407114 330664 407120 330676
rect 352064 330636 407120 330664
rect 352064 330624 352070 330636
rect 407114 330624 407120 330636
rect 407172 330624 407178 330676
rect 213914 330556 213920 330608
rect 213972 330596 213978 330608
rect 306926 330596 306932 330608
rect 213972 330568 306932 330596
rect 213972 330556 213978 330568
rect 306926 330556 306932 330568
rect 306984 330556 306990 330608
rect 327350 330556 327356 330608
rect 327408 330556 327414 330608
rect 334342 330556 334348 330608
rect 334400 330556 334406 330608
rect 373350 330556 373356 330608
rect 373408 330596 373414 330608
rect 498194 330596 498200 330608
rect 373408 330568 498200 330596
rect 373408 330556 373414 330568
rect 498194 330556 498200 330568
rect 498252 330556 498258 330608
rect 103514 330488 103520 330540
rect 103572 330528 103578 330540
rect 103572 330500 278912 330528
rect 103572 330488 103578 330500
rect 273438 330420 273444 330472
rect 273496 330460 273502 330472
rect 274082 330460 274088 330472
rect 273496 330432 274088 330460
rect 273496 330420 273502 330432
rect 274082 330420 274088 330432
rect 274140 330420 274146 330472
rect 274818 330420 274824 330472
rect 274876 330460 274882 330472
rect 275462 330460 275468 330472
rect 274876 330432 275468 330460
rect 274876 330420 274882 330432
rect 275462 330420 275468 330432
rect 275520 330420 275526 330472
rect 277394 330420 277400 330472
rect 277452 330460 277458 330472
rect 278222 330460 278228 330472
rect 277452 330432 278228 330460
rect 277452 330420 277458 330432
rect 278222 330420 278228 330432
rect 278280 330420 278286 330472
rect 278884 330460 278912 330500
rect 278958 330488 278964 330540
rect 279016 330528 279022 330540
rect 279602 330528 279608 330540
rect 279016 330500 279608 330528
rect 279016 330488 279022 330500
rect 279602 330488 279608 330500
rect 279660 330488 279666 330540
rect 281626 330488 281632 330540
rect 281684 330528 281690 330540
rect 282362 330528 282368 330540
rect 281684 330500 282368 330528
rect 281684 330488 281690 330500
rect 282362 330488 282368 330500
rect 282420 330488 282426 330540
rect 282914 330488 282920 330540
rect 282972 330528 282978 330540
rect 283466 330528 283472 330540
rect 282972 330500 283472 330528
rect 282972 330488 282978 330500
rect 283466 330488 283472 330500
rect 283524 330488 283530 330540
rect 284386 330488 284392 330540
rect 284444 330528 284450 330540
rect 285398 330528 285404 330540
rect 284444 330500 285404 330528
rect 284444 330488 284450 330500
rect 285398 330488 285404 330500
rect 285456 330488 285462 330540
rect 285950 330488 285956 330540
rect 286008 330528 286014 330540
rect 286502 330528 286508 330540
rect 286008 330500 286508 330528
rect 286008 330488 286014 330500
rect 286502 330488 286508 330500
rect 286560 330488 286566 330540
rect 287330 330488 287336 330540
rect 287388 330528 287394 330540
rect 288158 330528 288164 330540
rect 287388 330500 288164 330528
rect 287388 330488 287394 330500
rect 288158 330488 288164 330500
rect 288216 330488 288222 330540
rect 288710 330488 288716 330540
rect 288768 330528 288774 330540
rect 289262 330528 289268 330540
rect 288768 330500 289268 330528
rect 288768 330488 288774 330500
rect 289262 330488 289268 330500
rect 289320 330488 289326 330540
rect 291562 330488 291568 330540
rect 291620 330528 291626 330540
rect 292298 330528 292304 330540
rect 291620 330500 292304 330528
rect 291620 330488 291626 330500
rect 292298 330488 292304 330500
rect 292356 330488 292362 330540
rect 292666 330488 292672 330540
rect 292724 330528 292730 330540
rect 293678 330528 293684 330540
rect 292724 330500 293684 330528
rect 292724 330488 292730 330500
rect 293678 330488 293684 330500
rect 293736 330488 293742 330540
rect 296990 330488 296996 330540
rect 297048 330528 297054 330540
rect 297818 330528 297824 330540
rect 297048 330500 297824 330528
rect 297048 330488 297054 330500
rect 297818 330488 297824 330500
rect 297876 330488 297882 330540
rect 298186 330488 298192 330540
rect 298244 330528 298250 330540
rect 298922 330528 298928 330540
rect 298244 330500 298928 330528
rect 298244 330488 298250 330500
rect 298922 330488 298928 330500
rect 298980 330488 298986 330540
rect 301130 330488 301136 330540
rect 301188 330528 301194 330540
rect 301958 330528 301964 330540
rect 301188 330500 301964 330528
rect 301188 330488 301194 330500
rect 301958 330488 301964 330500
rect 302016 330488 302022 330540
rect 313642 330488 313648 330540
rect 313700 330528 313706 330540
rect 314102 330528 314108 330540
rect 313700 330500 314108 330528
rect 313700 330488 313706 330500
rect 314102 330488 314108 330500
rect 314160 330488 314166 330540
rect 317690 330488 317696 330540
rect 317748 330528 317754 330540
rect 318242 330528 318248 330540
rect 317748 330500 318248 330528
rect 317748 330488 317754 330500
rect 318242 330488 318248 330500
rect 318300 330488 318306 330540
rect 321646 330488 321652 330540
rect 321704 330528 321710 330540
rect 322382 330528 322388 330540
rect 321704 330500 322388 330528
rect 321704 330488 321710 330500
rect 322382 330488 322388 330500
rect 322440 330488 322446 330540
rect 323210 330488 323216 330540
rect 323268 330528 323274 330540
rect 324038 330528 324044 330540
rect 323268 330500 324044 330528
rect 323268 330488 323274 330500
rect 324038 330488 324044 330500
rect 324096 330488 324102 330540
rect 324406 330488 324412 330540
rect 324464 330528 324470 330540
rect 325142 330528 325148 330540
rect 324464 330500 325148 330528
rect 324464 330488 324470 330500
rect 325142 330488 325148 330500
rect 325200 330488 325206 330540
rect 327166 330488 327172 330540
rect 327224 330528 327230 330540
rect 328178 330528 328184 330540
rect 327224 330500 328184 330528
rect 327224 330488 327230 330500
rect 328178 330488 328184 330500
rect 328236 330488 328242 330540
rect 328730 330488 328736 330540
rect 328788 330528 328794 330540
rect 329558 330528 329564 330540
rect 328788 330500 329564 330528
rect 328788 330488 328794 330500
rect 329558 330488 329564 330500
rect 329616 330488 329622 330540
rect 331306 330488 331312 330540
rect 331364 330528 331370 330540
rect 332318 330528 332324 330540
rect 331364 330500 332324 330528
rect 331364 330488 331370 330500
rect 332318 330488 332324 330500
rect 332376 330488 332382 330540
rect 332686 330488 332692 330540
rect 332744 330528 332750 330540
rect 333422 330528 333428 330540
rect 332744 330500 333428 330528
rect 332744 330488 332750 330500
rect 333422 330488 333428 330500
rect 333480 330488 333486 330540
rect 334250 330488 334256 330540
rect 334308 330528 334314 330540
rect 334802 330528 334808 330540
rect 334308 330500 334808 330528
rect 334308 330488 334314 330500
rect 334802 330488 334808 330500
rect 334860 330488 334866 330540
rect 335446 330488 335452 330540
rect 335504 330528 335510 330540
rect 336458 330528 336464 330540
rect 335504 330500 336464 330528
rect 335504 330488 335510 330500
rect 336458 330488 336464 330500
rect 336516 330488 336522 330540
rect 336826 330488 336832 330540
rect 336884 330528 336890 330540
rect 337286 330528 337292 330540
rect 336884 330500 337292 330528
rect 336884 330488 336890 330500
rect 337286 330488 337292 330500
rect 337344 330488 337350 330540
rect 338206 330488 338212 330540
rect 338264 330528 338270 330540
rect 338942 330528 338948 330540
rect 338264 330500 338948 330528
rect 338264 330488 338270 330500
rect 338942 330488 338948 330500
rect 339000 330488 339006 330540
rect 339494 330488 339500 330540
rect 339552 330528 339558 330540
rect 340598 330528 340604 330540
rect 339552 330500 340604 330528
rect 339552 330488 339558 330500
rect 340598 330488 340604 330500
rect 340656 330488 340662 330540
rect 360286 330488 360292 330540
rect 360344 330528 360350 330540
rect 361022 330528 361028 330540
rect 360344 330500 361028 330528
rect 360344 330488 360350 330500
rect 361022 330488 361028 330500
rect 361080 330488 361086 330540
rect 361574 330488 361580 330540
rect 361632 330528 361638 330540
rect 362678 330528 362684 330540
rect 361632 330500 362684 330528
rect 361632 330488 361638 330500
rect 362678 330488 362684 330500
rect 362736 330488 362742 330540
rect 363138 330488 363144 330540
rect 363196 330528 363202 330540
rect 364058 330528 364064 330540
rect 363196 330500 364064 330528
rect 363196 330488 363202 330500
rect 364058 330488 364064 330500
rect 364116 330488 364122 330540
rect 364518 330488 364524 330540
rect 364576 330528 364582 330540
rect 365162 330528 365168 330540
rect 364576 330500 365168 330528
rect 364576 330488 364582 330500
rect 365162 330488 365168 330500
rect 365220 330488 365226 330540
rect 365714 330488 365720 330540
rect 365772 330528 365778 330540
rect 366266 330528 366272 330540
rect 365772 330500 366272 330528
rect 365772 330488 365778 330500
rect 366266 330488 366272 330500
rect 366324 330488 366330 330540
rect 368474 330488 368480 330540
rect 368532 330528 368538 330540
rect 368750 330528 368756 330540
rect 368532 330500 368756 330528
rect 368532 330488 368538 330500
rect 368750 330488 368756 330500
rect 368808 330488 368814 330540
rect 389450 330488 389456 330540
rect 389508 330528 389514 330540
rect 390002 330528 390008 330540
rect 389508 330500 390008 330528
rect 389508 330488 389514 330500
rect 390002 330488 390008 330500
rect 390060 330488 390066 330540
rect 390830 330488 390836 330540
rect 390888 330528 390894 330540
rect 391658 330528 391664 330540
rect 390888 330500 391664 330528
rect 390888 330488 390894 330500
rect 391658 330488 391664 330500
rect 391716 330488 391722 330540
rect 391934 330488 391940 330540
rect 391992 330528 391998 330540
rect 392486 330528 392492 330540
rect 391992 330500 392492 330528
rect 391992 330488 391998 330500
rect 392486 330488 392492 330500
rect 392544 330488 392550 330540
rect 571978 330528 571984 330540
rect 393286 330500 571984 330528
rect 281258 330460 281264 330472
rect 278884 330432 281264 330460
rect 281258 330420 281264 330432
rect 281316 330420 281322 330472
rect 283006 330420 283012 330472
rect 283064 330460 283070 330472
rect 284018 330460 284024 330472
rect 283064 330432 284024 330460
rect 283064 330420 283070 330432
rect 284018 330420 284024 330432
rect 284076 330420 284082 330472
rect 285858 330420 285864 330472
rect 285916 330460 285922 330472
rect 286778 330460 286784 330472
rect 285916 330432 286784 330460
rect 285916 330420 285922 330432
rect 286778 330420 286784 330432
rect 286836 330420 286842 330472
rect 288618 330420 288624 330472
rect 288676 330460 288682 330472
rect 289538 330460 289544 330472
rect 288676 330432 289544 330460
rect 288676 330420 288682 330432
rect 289538 330420 289544 330432
rect 289596 330420 289602 330472
rect 292850 330420 292856 330472
rect 292908 330460 292914 330472
rect 293402 330460 293408 330472
rect 292908 330432 293408 330460
rect 292908 330420 292914 330432
rect 293402 330420 293408 330432
rect 293460 330420 293466 330472
rect 298278 330420 298284 330472
rect 298336 330460 298342 330472
rect 299198 330460 299204 330472
rect 298336 330432 299204 330460
rect 298336 330420 298342 330432
rect 299198 330420 299204 330432
rect 299256 330420 299262 330472
rect 313458 330420 313464 330472
rect 313516 330460 313522 330472
rect 314378 330460 314384 330472
rect 313516 330432 314384 330460
rect 313516 330420 313522 330432
rect 314378 330420 314384 330432
rect 314436 330420 314442 330472
rect 315022 330420 315028 330472
rect 315080 330460 315086 330472
rect 315482 330460 315488 330472
rect 315080 330432 315488 330460
rect 315080 330420 315086 330432
rect 315482 330420 315488 330432
rect 315540 330420 315546 330472
rect 317506 330420 317512 330472
rect 317564 330460 317570 330472
rect 318518 330460 318524 330472
rect 317564 330432 318524 330460
rect 317564 330420 317570 330432
rect 318518 330420 318524 330432
rect 318576 330420 318582 330472
rect 324498 330420 324504 330472
rect 324556 330460 324562 330472
rect 325418 330460 325424 330472
rect 324556 330432 325424 330460
rect 324556 330420 324562 330432
rect 325418 330420 325424 330432
rect 325476 330420 325482 330472
rect 327442 330420 327448 330472
rect 327500 330460 327506 330472
rect 327902 330460 327908 330472
rect 327500 330432 327908 330460
rect 327500 330420 327506 330432
rect 327902 330420 327908 330432
rect 327960 330420 327966 330472
rect 328454 330420 328460 330472
rect 328512 330460 328518 330472
rect 329006 330460 329012 330472
rect 328512 330432 329012 330460
rect 328512 330420 328518 330432
rect 329006 330420 329012 330432
rect 329064 330420 329070 330472
rect 332870 330420 332876 330472
rect 332928 330460 332934 330472
rect 333146 330460 333152 330472
rect 332928 330432 333152 330460
rect 332928 330420 332934 330432
rect 333146 330420 333152 330432
rect 333204 330420 333210 330472
rect 333974 330420 333980 330472
rect 334032 330460 334038 330472
rect 335078 330460 335084 330472
rect 334032 330432 335084 330460
rect 334032 330420 334038 330432
rect 335078 330420 335084 330432
rect 335136 330420 335142 330472
rect 336918 330420 336924 330472
rect 336976 330460 336982 330472
rect 337562 330460 337568 330472
rect 336976 330432 337568 330460
rect 336976 330420 336982 330432
rect 337562 330420 337568 330432
rect 337620 330420 337626 330472
rect 338298 330420 338304 330472
rect 338356 330460 338362 330472
rect 339218 330460 339224 330472
rect 338356 330432 339224 330460
rect 338356 330420 338362 330432
rect 339218 330420 339224 330432
rect 339276 330420 339282 330472
rect 360194 330420 360200 330472
rect 360252 330460 360258 330472
rect 361298 330460 361304 330472
rect 360252 330432 361304 330460
rect 360252 330420 360258 330432
rect 361298 330420 361304 330432
rect 361356 330420 361362 330472
rect 364426 330420 364432 330472
rect 364484 330460 364490 330472
rect 365438 330460 365444 330472
rect 364484 330432 365444 330460
rect 364484 330420 364490 330432
rect 365438 330420 365444 330432
rect 365496 330420 365502 330472
rect 365806 330420 365812 330472
rect 365864 330460 365870 330472
rect 366818 330460 366824 330472
rect 365864 330432 366824 330460
rect 365864 330420 365870 330432
rect 366818 330420 366824 330432
rect 366876 330420 366882 330472
rect 368566 330420 368572 330472
rect 368624 330460 368630 330472
rect 369578 330460 369584 330472
rect 368624 330432 369584 330460
rect 368624 330420 368630 330432
rect 369578 330420 369584 330432
rect 369636 330420 369642 330472
rect 392026 330420 392032 330472
rect 392084 330460 392090 330472
rect 392762 330460 392768 330472
rect 392084 330432 392768 330460
rect 392084 330420 392090 330432
rect 392762 330420 392768 330432
rect 392820 330420 392826 330472
rect 273346 330352 273352 330404
rect 273404 330392 273410 330404
rect 274358 330392 274364 330404
rect 273404 330364 274364 330392
rect 273404 330352 273410 330364
rect 274358 330352 274364 330364
rect 274416 330352 274422 330404
rect 274726 330352 274732 330404
rect 274784 330392 274790 330404
rect 275738 330392 275744 330404
rect 274784 330364 275744 330392
rect 274784 330352 274790 330364
rect 275738 330352 275744 330364
rect 275796 330352 275802 330404
rect 283190 330352 283196 330404
rect 283248 330392 283254 330404
rect 283742 330392 283748 330404
rect 283248 330364 283748 330392
rect 283248 330352 283254 330364
rect 283742 330352 283748 330364
rect 283800 330352 283806 330404
rect 299842 330352 299848 330404
rect 299900 330392 299906 330404
rect 300578 330392 300584 330404
rect 299900 330364 300584 330392
rect 299900 330352 299906 330364
rect 300578 330352 300584 330364
rect 300636 330352 300642 330404
rect 390554 330352 390560 330404
rect 390612 330392 390618 330404
rect 393286 330392 393314 330500
rect 571978 330488 571984 330500
rect 572036 330488 572042 330540
rect 390612 330364 393314 330392
rect 390612 330352 390618 330364
rect 299658 330284 299664 330336
rect 299716 330324 299722 330336
rect 300302 330324 300308 330336
rect 299716 330296 300308 330324
rect 299716 330284 299722 330296
rect 300302 330284 300308 330296
rect 300360 330284 300366 330336
rect 332778 330148 332784 330200
rect 332836 330188 332842 330200
rect 333698 330188 333704 330200
rect 332836 330160 333704 330188
rect 332836 330148 332842 330160
rect 333698 330148 333704 330160
rect 333756 330148 333762 330200
rect 277670 329808 277676 329860
rect 277728 329848 277734 329860
rect 277946 329848 277952 329860
rect 277728 329820 277952 329848
rect 277728 329808 277734 329820
rect 277946 329808 277952 329820
rect 278004 329808 278010 329860
rect 323118 329740 323124 329792
rect 323176 329780 323182 329792
rect 323762 329780 323768 329792
rect 323176 329752 323768 329780
rect 323176 329740 323182 329752
rect 323762 329740 323768 329752
rect 323820 329740 323826 329792
rect 389266 329400 389272 329452
rect 389324 329440 389330 329452
rect 390278 329440 390284 329452
rect 389324 329412 390284 329440
rect 389324 329400 389330 329412
rect 390278 329400 390284 329412
rect 390336 329400 390342 329452
rect 277578 329264 277584 329316
rect 277636 329304 277642 329316
rect 278498 329304 278504 329316
rect 277636 329276 278504 329304
rect 277636 329264 277642 329276
rect 278498 329264 278504 329276
rect 278556 329264 278562 329316
rect 360562 329196 360568 329248
rect 360620 329236 360626 329248
rect 426434 329236 426440 329248
rect 360620 329208 426440 329236
rect 360620 329196 360626 329208
rect 426434 329196 426440 329208
rect 426492 329196 426498 329248
rect 224954 329128 224960 329180
rect 225012 329168 225018 329180
rect 309594 329168 309600 329180
rect 225012 329140 309600 329168
rect 225012 329128 225018 329140
rect 309594 329128 309600 329140
rect 309652 329128 309658 329180
rect 375926 329128 375932 329180
rect 375984 329168 375990 329180
rect 507854 329168 507860 329180
rect 375984 329140 507860 329168
rect 375984 329128 375990 329140
rect 507854 329128 507860 329140
rect 507912 329128 507918 329180
rect 149054 329060 149060 329112
rect 149112 329100 149118 329112
rect 291746 329100 291752 329112
rect 149112 329072 291752 329100
rect 149112 329060 149118 329072
rect 291746 329060 291752 329072
rect 291804 329060 291810 329112
rect 384390 329060 384396 329112
rect 384448 329100 384454 329112
rect 545114 329100 545120 329112
rect 384448 329072 545120 329100
rect 384448 329060 384454 329072
rect 545114 329060 545120 329072
rect 545172 329060 545178 329112
rect 364242 328516 364248 328568
rect 364300 328556 364306 328568
rect 364702 328556 364708 328568
rect 364300 328528 364708 328556
rect 364300 328516 364306 328528
rect 364702 328516 364708 328528
rect 364760 328516 364766 328568
rect 311986 328312 311992 328364
rect 312044 328352 312050 328364
rect 312998 328352 313004 328364
rect 312044 328324 313004 328352
rect 312044 328312 312050 328324
rect 312998 328312 313004 328324
rect 313056 328312 313062 328364
rect 367186 328176 367192 328228
rect 367244 328216 367250 328228
rect 367922 328216 367928 328228
rect 367244 328188 367928 328216
rect 367244 328176 367250 328188
rect 367922 328176 367928 328188
rect 367980 328176 367986 328228
rect 320450 328040 320456 328092
rect 320508 328080 320514 328092
rect 321278 328080 321284 328092
rect 320508 328052 321284 328080
rect 320508 328040 320514 328052
rect 321278 328040 321284 328052
rect 321336 328040 321342 328092
rect 339586 328040 339592 328092
rect 339644 328080 339650 328092
rect 340322 328080 340328 328092
rect 339644 328052 340328 328080
rect 339644 328040 339650 328052
rect 340322 328040 340328 328052
rect 340380 328040 340386 328092
rect 361666 327904 361672 327956
rect 361724 327944 361730 327956
rect 362402 327944 362408 327956
rect 361724 327916 362408 327944
rect 361724 327904 361730 327916
rect 362402 327904 362408 327916
rect 362460 327904 362466 327956
rect 189074 327836 189080 327888
rect 189132 327876 189138 327888
rect 300854 327876 300860 327888
rect 189132 327848 300860 327876
rect 189132 327836 189138 327848
rect 300854 327836 300860 327848
rect 300912 327836 300918 327888
rect 161474 327768 161480 327820
rect 161532 327808 161538 327820
rect 294782 327808 294788 327820
rect 161532 327780 294788 327808
rect 161532 327768 161538 327780
rect 294782 327768 294788 327780
rect 294840 327768 294846 327820
rect 363690 327768 363696 327820
rect 363748 327808 363754 327820
rect 448514 327808 448520 327820
rect 363748 327780 448520 327808
rect 363748 327768 363754 327780
rect 448514 327768 448520 327780
rect 448572 327768 448578 327820
rect 85574 327700 85580 327752
rect 85632 327740 85638 327752
rect 277118 327740 277124 327752
rect 85632 327712 277124 327740
rect 85632 327700 85638 327712
rect 277118 327700 277124 327712
rect 277176 327700 277182 327752
rect 314746 327700 314752 327752
rect 314804 327740 314810 327752
rect 315758 327740 315764 327752
rect 314804 327712 315764 327740
rect 314804 327700 314810 327712
rect 315758 327700 315764 327712
rect 315816 327700 315822 327752
rect 376478 327700 376484 327752
rect 376536 327740 376542 327752
rect 511994 327740 512000 327752
rect 376536 327712 512000 327740
rect 376536 327700 376542 327712
rect 511994 327700 512000 327712
rect 512052 327700 512058 327752
rect 291286 327020 291292 327072
rect 291344 327060 291350 327072
rect 292022 327060 292028 327072
rect 291344 327032 292028 327060
rect 291344 327020 291350 327032
rect 292022 327020 292028 327032
rect 292080 327020 292086 327072
rect 319070 326884 319076 326936
rect 319128 326924 319134 326936
rect 319898 326924 319904 326936
rect 319128 326896 319904 326924
rect 319128 326884 319134 326896
rect 319898 326884 319904 326896
rect 319956 326884 319962 326936
rect 269390 326680 269396 326732
rect 269448 326720 269454 326732
rect 269574 326720 269580 326732
rect 269448 326692 269580 326720
rect 269448 326680 269454 326692
rect 269574 326680 269580 326692
rect 269632 326680 269638 326732
rect 363046 326612 363052 326664
rect 363104 326652 363110 326664
rect 363506 326652 363512 326664
rect 363104 326624 363512 326652
rect 363104 326612 363110 326624
rect 363506 326612 363512 326624
rect 363564 326612 363570 326664
rect 263778 326544 263784 326596
rect 263836 326584 263842 326596
rect 264054 326584 264060 326596
rect 263836 326556 264060 326584
rect 263836 326544 263842 326556
rect 264054 326544 264060 326556
rect 264112 326544 264118 326596
rect 269298 326544 269304 326596
rect 269356 326584 269362 326596
rect 269482 326584 269488 326596
rect 269356 326556 269488 326584
rect 269356 326544 269362 326556
rect 269482 326544 269488 326556
rect 269540 326544 269546 326596
rect 320266 326544 320272 326596
rect 320324 326584 320330 326596
rect 321002 326584 321008 326596
rect 320324 326556 321008 326584
rect 320324 326544 320330 326556
rect 321002 326544 321008 326556
rect 321060 326544 321066 326596
rect 201494 326476 201500 326528
rect 201552 326516 201558 326528
rect 303614 326516 303620 326528
rect 201552 326488 303620 326516
rect 201552 326476 201558 326488
rect 303614 326476 303620 326488
rect 303672 326476 303678 326528
rect 382366 326476 382372 326528
rect 382424 326516 382430 326528
rect 383378 326516 383384 326528
rect 382424 326488 383384 326516
rect 382424 326476 382430 326488
rect 383378 326476 383384 326488
rect 383436 326476 383442 326528
rect 385310 326476 385316 326528
rect 385368 326516 385374 326528
rect 385494 326516 385500 326528
rect 385368 326488 385500 326516
rect 385368 326476 385374 326488
rect 385494 326476 385500 326488
rect 385552 326476 385558 326528
rect 182174 326408 182180 326460
rect 182232 326448 182238 326460
rect 299474 326448 299480 326460
rect 182232 326420 299480 326448
rect 182232 326408 182238 326420
rect 299474 326408 299480 326420
rect 299532 326408 299538 326460
rect 302326 326408 302332 326460
rect 302384 326448 302390 326460
rect 303338 326448 303344 326460
rect 302384 326420 303344 326448
rect 302384 326408 302390 326420
rect 303338 326408 303344 326420
rect 303396 326408 303402 326460
rect 303982 326408 303988 326460
rect 304040 326448 304046 326460
rect 304442 326448 304448 326460
rect 304040 326420 304448 326448
rect 304040 326408 304046 326420
rect 304442 326408 304448 326420
rect 304500 326408 304506 326460
rect 305178 326408 305184 326460
rect 305236 326448 305242 326460
rect 306098 326448 306104 326460
rect 305236 326420 306104 326448
rect 305236 326408 305242 326420
rect 306098 326408 306104 326420
rect 306156 326408 306162 326460
rect 309318 326408 309324 326460
rect 309376 326448 309382 326460
rect 310238 326448 310244 326460
rect 309376 326420 310244 326448
rect 309376 326408 309382 326420
rect 310238 326408 310244 326420
rect 310296 326408 310302 326460
rect 345198 326408 345204 326460
rect 345256 326448 345262 326460
rect 346118 326448 346124 326460
rect 345256 326420 346124 326448
rect 345256 326408 345262 326420
rect 346118 326408 346124 326420
rect 346176 326408 346182 326460
rect 346394 326408 346400 326460
rect 346452 326448 346458 326460
rect 347498 326448 347504 326460
rect 346452 326420 347504 326448
rect 346452 326408 346458 326420
rect 347498 326408 347504 326420
rect 347556 326408 347562 326460
rect 347958 326408 347964 326460
rect 348016 326448 348022 326460
rect 348142 326448 348148 326460
rect 348016 326420 348148 326448
rect 348016 326408 348022 326420
rect 348142 326408 348148 326420
rect 348200 326408 348206 326460
rect 350718 326408 350724 326460
rect 350776 326448 350782 326460
rect 350994 326448 351000 326460
rect 350776 326420 351000 326448
rect 350776 326408 350782 326420
rect 350994 326408 351000 326420
rect 351052 326408 351058 326460
rect 353386 326408 353392 326460
rect 353444 326448 353450 326460
rect 354398 326448 354404 326460
rect 353444 326420 354404 326448
rect 353444 326408 353450 326420
rect 354398 326408 354404 326420
rect 354456 326408 354462 326460
rect 354766 326408 354772 326460
rect 354824 326448 354830 326460
rect 355502 326448 355508 326460
rect 354824 326420 355508 326448
rect 354824 326408 354830 326420
rect 355502 326408 355508 326420
rect 355560 326408 355566 326460
rect 357526 326408 357532 326460
rect 357584 326448 357590 326460
rect 358262 326448 358268 326460
rect 357584 326420 358268 326448
rect 357584 326408 357590 326420
rect 358262 326408 358268 326420
rect 358320 326408 358326 326460
rect 358906 326408 358912 326460
rect 358964 326448 358970 326460
rect 359918 326448 359924 326460
rect 358964 326420 359924 326448
rect 358964 326408 358970 326420
rect 359918 326408 359924 326420
rect 359976 326408 359982 326460
rect 364886 326408 364892 326460
rect 364944 326448 364950 326460
rect 462314 326448 462320 326460
rect 364944 326420 462320 326448
rect 364944 326408 364950 326420
rect 462314 326408 462320 326420
rect 462372 326408 462378 326460
rect 53834 326340 53840 326392
rect 53892 326380 53898 326392
rect 53892 326352 253934 326380
rect 53892 326340 53898 326352
rect 253906 326312 253934 326352
rect 256786 326340 256792 326392
rect 256844 326380 256850 326392
rect 257522 326380 257528 326392
rect 256844 326352 257528 326380
rect 256844 326340 256850 326352
rect 257522 326340 257528 326352
rect 257580 326340 257586 326392
rect 258166 326340 258172 326392
rect 258224 326380 258230 326392
rect 258902 326380 258908 326392
rect 258224 326352 258908 326380
rect 258224 326340 258230 326352
rect 258902 326340 258908 326352
rect 258960 326340 258966 326392
rect 259638 326340 259644 326392
rect 259696 326380 259702 326392
rect 260282 326380 260288 326392
rect 259696 326352 260288 326380
rect 259696 326340 259702 326352
rect 260282 326340 260288 326352
rect 260340 326340 260346 326392
rect 261202 326340 261208 326392
rect 261260 326380 261266 326392
rect 261662 326380 261668 326392
rect 261260 326352 261668 326380
rect 261260 326340 261266 326352
rect 261662 326340 261668 326352
rect 261720 326340 261726 326392
rect 262306 326340 262312 326392
rect 262364 326380 262370 326392
rect 262766 326380 262772 326392
rect 262364 326352 262772 326380
rect 262364 326340 262370 326352
rect 262766 326340 262772 326352
rect 262824 326340 262830 326392
rect 264974 326340 264980 326392
rect 265032 326380 265038 326392
rect 265434 326380 265440 326392
rect 265032 326352 265440 326380
rect 265032 326340 265038 326352
rect 265434 326340 265440 326352
rect 265492 326340 265498 326392
rect 266446 326340 266452 326392
rect 266504 326380 266510 326392
rect 267458 326380 267464 326392
rect 266504 326352 267464 326380
rect 266504 326340 266510 326352
rect 267458 326340 267464 326352
rect 267516 326340 267522 326392
rect 267826 326340 267832 326392
rect 267884 326380 267890 326392
rect 268562 326380 268568 326392
rect 267884 326352 268568 326380
rect 267884 326340 267890 326352
rect 268562 326340 268568 326352
rect 268620 326340 268626 326392
rect 269482 326340 269488 326392
rect 269540 326380 269546 326392
rect 269942 326380 269948 326392
rect 269540 326352 269948 326380
rect 269540 326340 269546 326352
rect 269942 326340 269948 326352
rect 270000 326340 270006 326392
rect 270862 326340 270868 326392
rect 270920 326380 270926 326392
rect 271598 326380 271604 326392
rect 270920 326352 271604 326380
rect 270920 326340 270926 326352
rect 271598 326340 271604 326352
rect 271656 326340 271662 326392
rect 302602 326340 302608 326392
rect 302660 326380 302666 326392
rect 303062 326380 303068 326392
rect 302660 326352 303068 326380
rect 302660 326340 302666 326352
rect 303062 326340 303068 326352
rect 303120 326340 303126 326392
rect 303798 326340 303804 326392
rect 303856 326380 303862 326392
rect 304166 326380 304172 326392
rect 303856 326352 304172 326380
rect 303856 326340 303862 326352
rect 304166 326340 304172 326352
rect 304224 326340 304230 326392
rect 305270 326340 305276 326392
rect 305328 326380 305334 326392
rect 305822 326380 305828 326392
rect 305328 326352 305828 326380
rect 305328 326340 305334 326352
rect 305822 326340 305828 326352
rect 305880 326340 305886 326392
rect 306650 326340 306656 326392
rect 306708 326380 306714 326392
rect 307478 326380 307484 326392
rect 306708 326352 307484 326380
rect 306708 326340 306714 326352
rect 307478 326340 307484 326352
rect 307536 326340 307542 326392
rect 307846 326340 307852 326392
rect 307904 326380 307910 326392
rect 308306 326380 308312 326392
rect 307904 326352 308312 326380
rect 307904 326340 307910 326352
rect 308306 326340 308312 326352
rect 308364 326340 308370 326392
rect 309502 326340 309508 326392
rect 309560 326380 309566 326392
rect 309962 326380 309968 326392
rect 309560 326352 309968 326380
rect 309560 326340 309566 326352
rect 309962 326340 309968 326352
rect 310020 326340 310026 326392
rect 340966 326340 340972 326392
rect 341024 326380 341030 326392
rect 341702 326380 341708 326392
rect 341024 326352 341708 326380
rect 341024 326340 341030 326352
rect 341702 326340 341708 326352
rect 341760 326340 341766 326392
rect 342346 326340 342352 326392
rect 342404 326380 342410 326392
rect 343358 326380 343364 326392
rect 342404 326352 343364 326380
rect 342404 326340 342410 326352
rect 343358 326340 343364 326352
rect 343416 326340 343422 326392
rect 343634 326340 343640 326392
rect 343692 326380 343698 326392
rect 344738 326380 344744 326392
rect 343692 326352 344744 326380
rect 343692 326340 343698 326352
rect 344738 326340 344744 326352
rect 344796 326340 344802 326392
rect 345106 326340 345112 326392
rect 345164 326380 345170 326392
rect 345566 326380 345572 326392
rect 345164 326352 345572 326380
rect 345164 326340 345170 326352
rect 345566 326340 345572 326352
rect 345624 326340 345630 326392
rect 346486 326340 346492 326392
rect 346544 326380 346550 326392
rect 347222 326380 347228 326392
rect 346544 326352 347228 326380
rect 346544 326340 346550 326352
rect 347222 326340 347228 326352
rect 347280 326340 347286 326392
rect 347774 326340 347780 326392
rect 347832 326380 347838 326392
rect 348878 326380 348884 326392
rect 347832 326352 348884 326380
rect 347832 326340 347838 326352
rect 348878 326340 348884 326352
rect 348936 326340 348942 326392
rect 349154 326340 349160 326392
rect 349212 326380 349218 326392
rect 350258 326380 350264 326392
rect 349212 326352 350264 326380
rect 349212 326340 349218 326352
rect 350258 326340 350264 326352
rect 350316 326340 350322 326392
rect 350626 326340 350632 326392
rect 350684 326380 350690 326392
rect 351362 326380 351368 326392
rect 350684 326352 351368 326380
rect 350684 326340 350690 326352
rect 351362 326340 351368 326352
rect 351420 326340 351426 326392
rect 351914 326340 351920 326392
rect 351972 326380 351978 326392
rect 353018 326380 353024 326392
rect 351972 326352 353024 326380
rect 351972 326340 351978 326352
rect 353018 326340 353024 326352
rect 353076 326340 353082 326392
rect 353294 326340 353300 326392
rect 353352 326380 353358 326392
rect 353846 326380 353852 326392
rect 353352 326352 353852 326380
rect 353352 326340 353358 326352
rect 353846 326340 353852 326352
rect 353904 326340 353910 326392
rect 354950 326340 354956 326392
rect 355008 326380 355014 326392
rect 355226 326380 355232 326392
rect 355008 326352 355232 326380
rect 355008 326340 355014 326352
rect 355226 326340 355232 326352
rect 355284 326340 355290 326392
rect 356146 326340 356152 326392
rect 356204 326380 356210 326392
rect 357158 326380 357164 326392
rect 356204 326352 357164 326380
rect 356204 326340 356210 326352
rect 357158 326340 357164 326352
rect 357216 326340 357222 326392
rect 357434 326340 357440 326392
rect 357492 326380 357498 326392
rect 357986 326380 357992 326392
rect 357492 326352 357992 326380
rect 357492 326340 357498 326352
rect 357986 326340 357992 326352
rect 358044 326340 358050 326392
rect 358814 326340 358820 326392
rect 358872 326380 358878 326392
rect 359642 326380 359648 326392
rect 358872 326352 359648 326380
rect 358872 326340 358878 326352
rect 359642 326340 359648 326352
rect 359700 326340 359706 326392
rect 369854 326340 369860 326392
rect 369912 326380 369918 326392
rect 370406 326380 370412 326392
rect 369912 326352 370412 326380
rect 369912 326340 369918 326352
rect 370406 326340 370412 326352
rect 370464 326340 370470 326392
rect 371326 326340 371332 326392
rect 371384 326380 371390 326392
rect 372062 326380 372068 326392
rect 371384 326352 372068 326380
rect 371384 326340 371390 326352
rect 372062 326340 372068 326352
rect 372120 326340 372126 326392
rect 372890 326340 372896 326392
rect 372948 326380 372954 326392
rect 373442 326380 373448 326392
rect 372948 326352 373448 326380
rect 372948 326340 372954 326352
rect 373442 326340 373448 326352
rect 373500 326340 373506 326392
rect 374178 326340 374184 326392
rect 374236 326380 374242 326392
rect 374546 326380 374552 326392
rect 374236 326352 374552 326380
rect 374236 326340 374242 326352
rect 374546 326340 374552 326352
rect 374604 326340 374610 326392
rect 375374 326340 375380 326392
rect 375432 326380 375438 326392
rect 376294 326380 376300 326392
rect 375432 326352 376300 326380
rect 375432 326340 375438 326352
rect 376294 326340 376300 326352
rect 376352 326340 376358 326392
rect 378226 326340 378232 326392
rect 378284 326380 378290 326392
rect 378962 326380 378968 326392
rect 378284 326352 378968 326380
rect 378284 326340 378290 326352
rect 378962 326340 378968 326352
rect 379020 326340 379026 326392
rect 379514 326340 379520 326392
rect 379572 326380 379578 326392
rect 380342 326380 380348 326392
rect 379572 326352 380348 326380
rect 379572 326340 379578 326352
rect 380342 326340 380348 326352
rect 380400 326340 380406 326392
rect 381078 326340 381084 326392
rect 381136 326380 381142 326392
rect 381722 326380 381728 326392
rect 381136 326352 381728 326380
rect 381136 326340 381142 326352
rect 381722 326340 381728 326352
rect 381780 326340 381786 326392
rect 382458 326340 382464 326392
rect 382516 326380 382522 326392
rect 383102 326380 383108 326392
rect 382516 326352 383108 326380
rect 382516 326340 382522 326352
rect 383102 326340 383108 326352
rect 383160 326340 383166 326392
rect 383654 326340 383660 326392
rect 383712 326380 383718 326392
rect 384482 326380 384488 326392
rect 383712 326352 384488 326380
rect 383712 326340 383718 326352
rect 384482 326340 384488 326352
rect 384540 326340 384546 326392
rect 385034 326340 385040 326392
rect 385092 326380 385098 326392
rect 385862 326380 385868 326392
rect 385092 326352 385868 326380
rect 385092 326340 385098 326352
rect 385862 326340 385868 326352
rect 385920 326340 385926 326392
rect 386690 326340 386696 326392
rect 386748 326380 386754 326392
rect 387242 326380 387248 326392
rect 386748 326352 387248 326380
rect 386748 326340 386754 326352
rect 387242 326340 387248 326352
rect 387300 326340 387306 326392
rect 388070 326340 388076 326392
rect 388128 326380 388134 326392
rect 388898 326380 388904 326392
rect 388128 326352 388904 326380
rect 388128 326340 388134 326352
rect 388898 326340 388904 326352
rect 388956 326340 388962 326392
rect 525794 326380 525800 326392
rect 389146 326352 525800 326380
rect 253906 326284 268424 326312
rect 259546 326204 259552 326256
rect 259604 326244 259610 326256
rect 260558 326244 260564 326256
rect 259604 326216 260564 326244
rect 259604 326204 259610 326216
rect 260558 326204 260564 326216
rect 260616 326204 260622 326256
rect 260926 326204 260932 326256
rect 260984 326244 260990 326256
rect 261386 326244 261392 326256
rect 260984 326216 261392 326244
rect 260984 326204 260990 326216
rect 261386 326204 261392 326216
rect 261444 326204 261450 326256
rect 262398 326204 262404 326256
rect 262456 326244 262462 326256
rect 263318 326244 263324 326256
rect 262456 326216 263324 326244
rect 262456 326204 262462 326216
rect 263318 326204 263324 326216
rect 263376 326204 263382 326256
rect 263962 326204 263968 326256
rect 264020 326244 264026 326256
rect 264422 326244 264428 326256
rect 264020 326216 264428 326244
rect 264020 326204 264026 326216
rect 264422 326204 264428 326216
rect 264480 326204 264486 326256
rect 265158 326204 265164 326256
rect 265216 326244 265222 326256
rect 265802 326244 265808 326256
rect 265216 326216 265808 326244
rect 265216 326204 265222 326216
rect 265802 326204 265808 326216
rect 265860 326204 265866 326256
rect 267918 326204 267924 326256
rect 267976 326244 267982 326256
rect 268286 326244 268292 326256
rect 267976 326216 268292 326244
rect 267976 326204 267982 326216
rect 268286 326204 268292 326216
rect 268344 326204 268350 326256
rect 268396 326244 268424 326284
rect 269206 326272 269212 326324
rect 269264 326312 269270 326324
rect 270218 326312 270224 326324
rect 269264 326284 270224 326312
rect 269264 326272 269270 326284
rect 270218 326272 270224 326284
rect 270276 326272 270282 326324
rect 270770 326272 270776 326324
rect 270828 326312 270834 326324
rect 271322 326312 271328 326324
rect 270828 326284 271328 326312
rect 270828 326272 270834 326284
rect 271322 326272 271328 326284
rect 271380 326272 271386 326324
rect 303706 326272 303712 326324
rect 303764 326312 303770 326324
rect 304718 326312 304724 326324
rect 303764 326284 304724 326312
rect 303764 326272 303770 326284
rect 304718 326272 304724 326284
rect 304776 326272 304782 326324
rect 345014 326272 345020 326324
rect 345072 326312 345078 326324
rect 345842 326312 345848 326324
rect 345072 326284 345848 326312
rect 345072 326272 345078 326284
rect 345842 326272 345848 326284
rect 345900 326272 345906 326324
rect 357618 326272 357624 326324
rect 357676 326312 357682 326324
rect 358538 326312 358544 326324
rect 357676 326284 358544 326312
rect 357676 326272 357682 326284
rect 358538 326272 358544 326284
rect 358596 326272 358602 326324
rect 369946 326272 369952 326324
rect 370004 326312 370010 326324
rect 370958 326312 370964 326324
rect 370004 326284 370964 326312
rect 370004 326272 370010 326284
rect 370958 326272 370964 326284
rect 371016 326272 371022 326324
rect 372798 326272 372804 326324
rect 372856 326312 372862 326324
rect 373718 326312 373724 326324
rect 372856 326284 373724 326312
rect 372856 326272 372862 326284
rect 373718 326272 373724 326284
rect 373776 326272 373782 326324
rect 374270 326272 374276 326324
rect 374328 326312 374334 326324
rect 375098 326312 375104 326324
rect 374328 326284 375104 326312
rect 374328 326272 374334 326284
rect 375098 326272 375104 326284
rect 375156 326272 375162 326324
rect 378134 326272 378140 326324
rect 378192 326312 378198 326324
rect 379238 326312 379244 326324
rect 378192 326284 379244 326312
rect 378192 326272 378198 326284
rect 379238 326272 379244 326284
rect 379296 326272 379302 326324
rect 380986 326272 380992 326324
rect 381044 326312 381050 326324
rect 381998 326312 382004 326324
rect 381044 326284 382004 326312
rect 381044 326272 381050 326284
rect 381998 326272 382004 326284
rect 382056 326272 382062 326324
rect 382274 326272 382280 326324
rect 382332 326312 382338 326324
rect 382826 326312 382832 326324
rect 382332 326284 382832 326312
rect 382332 326272 382338 326284
rect 382826 326272 382832 326284
rect 382884 326272 382890 326324
rect 385126 326272 385132 326324
rect 385184 326312 385190 326324
rect 386138 326312 386144 326324
rect 385184 326284 386144 326312
rect 385184 326272 385190 326284
rect 386138 326272 386144 326284
rect 386196 326272 386202 326324
rect 386414 326272 386420 326324
rect 386472 326312 386478 326324
rect 386966 326312 386972 326324
rect 386472 326284 386972 326312
rect 386472 326272 386478 326284
rect 386966 326272 386972 326284
rect 387024 326272 387030 326324
rect 269666 326244 269672 326256
rect 268396 326216 269672 326244
rect 269666 326204 269672 326216
rect 269724 326204 269730 326256
rect 310606 326204 310612 326256
rect 310664 326244 310670 326256
rect 310790 326244 310796 326256
rect 310664 326216 310796 326244
rect 310664 326204 310670 326216
rect 310790 326204 310796 326216
rect 310848 326204 310854 326256
rect 310882 326204 310888 326256
rect 310940 326244 310946 326256
rect 311618 326244 311624 326256
rect 310940 326216 311624 326244
rect 310940 326204 310946 326216
rect 311618 326204 311624 326216
rect 311676 326204 311682 326256
rect 350810 326204 350816 326256
rect 350868 326244 350874 326256
rect 351638 326244 351644 326256
rect 350868 326216 351644 326244
rect 350868 326204 350874 326216
rect 351638 326204 351644 326216
rect 351696 326204 351702 326256
rect 376938 326204 376944 326256
rect 376996 326244 377002 326256
rect 377582 326244 377588 326256
rect 376996 326216 377588 326244
rect 376996 326204 377002 326216
rect 377582 326204 377588 326216
rect 377640 326204 377646 326256
rect 379790 326204 379796 326256
rect 379848 326244 379854 326256
rect 389146 326244 389174 326352
rect 525794 326340 525800 326352
rect 525852 326340 525858 326392
rect 379848 326216 389174 326244
rect 379848 326204 379854 326216
rect 265066 326136 265072 326188
rect 265124 326176 265130 326188
rect 266078 326176 266084 326188
rect 265124 326148 266084 326176
rect 265124 326136 265130 326148
rect 266078 326136 266084 326148
rect 266136 326136 266142 326188
rect 289906 326136 289912 326188
rect 289964 326176 289970 326188
rect 290642 326176 290648 326188
rect 289964 326148 290648 326176
rect 289964 326136 289970 326148
rect 290642 326136 290648 326148
rect 290700 326136 290706 326188
rect 376846 326136 376852 326188
rect 376904 326176 376910 326188
rect 377858 326176 377864 326188
rect 376904 326148 377864 326176
rect 376904 326136 376910 326148
rect 377858 326136 377864 326148
rect 377916 326136 377922 326188
rect 328546 325864 328552 325916
rect 328604 325904 328610 325916
rect 329282 325904 329288 325916
rect 328604 325876 329288 325904
rect 328604 325864 328610 325876
rect 329282 325864 329288 325876
rect 329340 325864 329346 325916
rect 368750 325864 368756 325916
rect 368808 325904 368814 325916
rect 369302 325904 369308 325916
rect 368808 325876 369308 325904
rect 368808 325864 368814 325876
rect 369302 325864 369308 325876
rect 369360 325864 369366 325916
rect 396810 325592 396816 325644
rect 396868 325632 396874 325644
rect 579890 325632 579896 325644
rect 396868 325604 579896 325632
rect 396868 325592 396874 325604
rect 579890 325592 579896 325604
rect 579948 325592 579954 325644
rect 266630 325320 266636 325372
rect 266688 325360 266694 325372
rect 267182 325360 267188 325372
rect 266688 325332 267188 325360
rect 266688 325320 266694 325332
rect 267182 325320 267188 325332
rect 267240 325320 267246 325372
rect 309226 325320 309232 325372
rect 309284 325360 309290 325372
rect 309686 325360 309692 325372
rect 309284 325332 309692 325360
rect 309284 325320 309290 325332
rect 309686 325320 309692 325332
rect 309744 325320 309750 325372
rect 231854 325048 231860 325100
rect 231912 325088 231918 325100
rect 311066 325088 311072 325100
rect 231912 325060 311072 325088
rect 231912 325048 231918 325060
rect 311066 325048 311072 325060
rect 311124 325048 311130 325100
rect 349798 325048 349804 325100
rect 349856 325088 349862 325100
rect 390554 325088 390560 325100
rect 349856 325060 390560 325088
rect 349856 325048 349862 325060
rect 390554 325048 390560 325060
rect 390612 325048 390618 325100
rect 164234 324980 164240 325032
rect 164292 325020 164298 325032
rect 295334 325020 295340 325032
rect 164292 324992 295340 325020
rect 164292 324980 164298 324992
rect 295334 324980 295340 324992
rect 295392 324980 295398 325032
rect 352466 324980 352472 325032
rect 352524 325020 352530 325032
rect 408494 325020 408500 325032
rect 352524 324992 408500 325020
rect 352524 324980 352530 324992
rect 408494 324980 408500 324992
rect 408552 324980 408558 325032
rect 46934 324912 46940 324964
rect 46992 324952 46998 324964
rect 268102 324952 268108 324964
rect 46992 324924 268108 324952
rect 46992 324912 46998 324924
rect 268102 324912 268108 324924
rect 268160 324912 268166 324964
rect 377214 324912 377220 324964
rect 377272 324952 377278 324964
rect 513374 324952 513380 324964
rect 377272 324924 513380 324952
rect 377272 324912 377278 324924
rect 513374 324912 513380 324924
rect 513432 324912 513438 324964
rect 386506 324640 386512 324692
rect 386564 324680 386570 324692
rect 387518 324680 387524 324692
rect 386564 324652 387524 324680
rect 386564 324640 386570 324652
rect 387518 324640 387524 324652
rect 387576 324640 387582 324692
rect 261110 324504 261116 324556
rect 261168 324544 261174 324556
rect 261938 324544 261944 324556
rect 261168 324516 261944 324544
rect 261168 324504 261174 324516
rect 261938 324504 261944 324516
rect 261996 324504 262002 324556
rect 343726 324368 343732 324420
rect 343784 324408 343790 324420
rect 344462 324408 344468 324420
rect 343784 324380 344468 324408
rect 343784 324368 343790 324380
rect 344462 324368 344468 324380
rect 344520 324368 344526 324420
rect 387794 324300 387800 324352
rect 387852 324340 387858 324352
rect 388622 324340 388628 324352
rect 387852 324312 388628 324340
rect 387852 324300 387858 324312
rect 388622 324300 388628 324312
rect 388680 324300 388686 324352
rect 310606 324232 310612 324284
rect 310664 324272 310670 324284
rect 311342 324272 311348 324284
rect 310664 324244 311348 324272
rect 310664 324232 310670 324244
rect 311342 324232 311348 324244
rect 311400 324232 311406 324284
rect 380894 324096 380900 324148
rect 380952 324136 380958 324148
rect 381262 324136 381268 324148
rect 380952 324108 381268 324136
rect 380952 324096 380958 324108
rect 381262 324096 381268 324108
rect 381320 324096 381326 324148
rect 238754 323756 238760 323808
rect 238812 323796 238818 323808
rect 309870 323796 309876 323808
rect 238812 323768 309876 323796
rect 238812 323756 238818 323768
rect 309870 323756 309876 323768
rect 309928 323756 309934 323808
rect 171134 323688 171140 323740
rect 171192 323728 171198 323740
rect 296254 323728 296260 323740
rect 171192 323700 296260 323728
rect 171192 323688 171198 323700
rect 296254 323688 296260 323700
rect 296312 323688 296318 323740
rect 306466 323688 306472 323740
rect 306524 323728 306530 323740
rect 307202 323728 307208 323740
rect 306524 323700 307208 323728
rect 306524 323688 306530 323700
rect 307202 323688 307208 323700
rect 307260 323688 307266 323740
rect 353662 323688 353668 323740
rect 353720 323728 353726 323740
rect 412634 323728 412640 323740
rect 353720 323700 412640 323728
rect 353720 323688 353726 323700
rect 412634 323688 412640 323700
rect 412692 323688 412698 323740
rect 155954 323620 155960 323672
rect 156012 323660 156018 323672
rect 292850 323660 292856 323672
rect 156012 323632 292856 323660
rect 156012 323620 156018 323632
rect 292850 323620 292856 323632
rect 292908 323620 292914 323672
rect 374822 323620 374828 323672
rect 374880 323660 374886 323672
rect 505094 323660 505100 323672
rect 374880 323632 505100 323660
rect 374880 323620 374886 323632
rect 505094 323620 505100 323632
rect 505152 323620 505158 323672
rect 25498 323552 25504 323604
rect 25556 323592 25562 323604
rect 262490 323592 262496 323604
rect 25556 323564 262496 323592
rect 25556 323552 25562 323564
rect 262490 323552 262496 323564
rect 262548 323552 262554 323604
rect 342438 323552 342444 323604
rect 342496 323592 342502 323604
rect 343082 323592 343088 323604
rect 342496 323564 343088 323592
rect 342496 323552 342502 323564
rect 343082 323552 343088 323564
rect 343140 323552 343146 323604
rect 359550 323552 359556 323604
rect 359608 323592 359614 323604
rect 373994 323592 374000 323604
rect 359608 323564 374000 323592
rect 359608 323552 359614 323564
rect 373994 323552 374000 323564
rect 374052 323552 374058 323604
rect 380066 323552 380072 323604
rect 380124 323592 380130 323604
rect 527174 323592 527180 323604
rect 380124 323564 527180 323592
rect 380124 323552 380130 323564
rect 527174 323552 527180 323564
rect 527232 323552 527238 323604
rect 387978 323212 387984 323264
rect 388036 323252 388042 323264
rect 388346 323252 388352 323264
rect 388036 323224 388352 323252
rect 388036 323212 388042 323224
rect 388346 323212 388352 323224
rect 388404 323212 388410 323264
rect 356330 323144 356336 323196
rect 356388 323184 356394 323196
rect 356882 323184 356888 323196
rect 356388 323156 356888 323184
rect 356388 323144 356394 323156
rect 356882 323144 356888 323156
rect 356940 323144 356946 323196
rect 354674 322736 354680 322788
rect 354732 322776 354738 322788
rect 355778 322776 355784 322788
rect 354732 322748 355784 322776
rect 354732 322736 354738 322748
rect 355778 322736 355784 322748
rect 355836 322736 355842 322788
rect 242986 322396 242992 322448
rect 243044 322436 243050 322448
rect 313550 322436 313556 322448
rect 243044 322408 313556 322436
rect 243044 322396 243050 322408
rect 313550 322396 313556 322408
rect 313608 322396 313614 322448
rect 175274 322328 175280 322380
rect 175332 322368 175338 322380
rect 296990 322368 296996 322380
rect 175332 322340 296996 322368
rect 175332 322328 175338 322340
rect 296990 322328 296996 322340
rect 297048 322328 297054 322380
rect 349246 322328 349252 322380
rect 349304 322368 349310 322380
rect 394694 322368 394700 322380
rect 349304 322340 394700 322368
rect 349304 322328 349310 322340
rect 394694 322328 394700 322340
rect 394752 322328 394758 322380
rect 142154 322260 142160 322312
rect 142212 322300 142218 322312
rect 289998 322300 290004 322312
rect 142212 322272 290004 322300
rect 142212 322260 142218 322272
rect 289998 322260 290004 322272
rect 290056 322260 290062 322312
rect 366542 322260 366548 322312
rect 366600 322300 366606 322312
rect 469214 322300 469220 322312
rect 366600 322272 469220 322300
rect 366600 322260 366606 322272
rect 469214 322260 469220 322272
rect 469272 322260 469278 322312
rect 34514 322192 34520 322244
rect 34572 322232 34578 322244
rect 265342 322232 265348 322244
rect 34572 322204 265348 322232
rect 34572 322192 34578 322204
rect 265342 322192 265348 322204
rect 265400 322192 265406 322244
rect 378502 322192 378508 322244
rect 378560 322232 378566 322244
rect 518894 322232 518900 322244
rect 378560 322204 518900 322232
rect 378560 322192 378566 322204
rect 518894 322192 518900 322204
rect 518952 322192 518958 322244
rect 346578 321648 346584 321700
rect 346636 321688 346642 321700
rect 346762 321688 346768 321700
rect 346636 321660 346768 321688
rect 346636 321648 346642 321660
rect 346762 321648 346768 321660
rect 346820 321648 346826 321700
rect 259730 321308 259736 321360
rect 259788 321348 259794 321360
rect 259914 321348 259920 321360
rect 259788 321320 259920 321348
rect 259788 321308 259794 321320
rect 259914 321308 259920 321320
rect 259972 321308 259978 321360
rect 249794 320968 249800 321020
rect 249852 321008 249858 321020
rect 314930 321008 314936 321020
rect 249852 320980 314936 321008
rect 249852 320968 249858 320980
rect 314930 320968 314936 320980
rect 314988 320968 314994 321020
rect 350902 320968 350908 321020
rect 350960 321008 350966 321020
rect 401594 321008 401600 321020
rect 350960 320980 401600 321008
rect 350960 320968 350966 320980
rect 401594 320968 401600 320980
rect 401652 320968 401658 321020
rect 178034 320900 178040 320952
rect 178092 320940 178098 320952
rect 297542 320940 297548 320952
rect 178092 320912 297548 320940
rect 178092 320900 178098 320912
rect 297542 320900 297548 320912
rect 297600 320900 297606 320952
rect 378226 320900 378232 320952
rect 378284 320940 378290 320952
rect 523034 320940 523040 320952
rect 378284 320912 523040 320940
rect 378284 320900 378290 320912
rect 523034 320900 523040 320912
rect 523092 320900 523098 320952
rect 131114 320832 131120 320884
rect 131172 320872 131178 320884
rect 286318 320872 286324 320884
rect 131172 320844 286324 320872
rect 131172 320832 131178 320844
rect 286318 320832 286324 320844
rect 286376 320832 286382 320884
rect 287054 320832 287060 320884
rect 287112 320872 287118 320884
rect 287238 320872 287244 320884
rect 287112 320844 287244 320872
rect 287112 320832 287118 320844
rect 287238 320832 287244 320844
rect 287296 320832 287302 320884
rect 389174 320832 389180 320884
rect 389232 320872 389238 320884
rect 565814 320872 565820 320884
rect 389232 320844 565820 320872
rect 389232 320832 389238 320844
rect 565814 320832 565820 320844
rect 565872 320832 565878 320884
rect 3510 320084 3516 320136
rect 3568 320124 3574 320136
rect 233970 320124 233976 320136
rect 3568 320096 233976 320124
rect 3568 320084 3574 320096
rect 233970 320084 233976 320096
rect 234028 320084 234034 320136
rect 252554 319540 252560 319592
rect 252612 319580 252618 319592
rect 305730 319580 305736 319592
rect 252612 319552 305736 319580
rect 252612 319540 252618 319552
rect 305730 319540 305736 319552
rect 305788 319540 305794 319592
rect 350810 319540 350816 319592
rect 350868 319580 350874 319592
rect 405734 319580 405740 319592
rect 350868 319552 405740 319580
rect 350868 319540 350874 319552
rect 405734 319540 405740 319552
rect 405792 319540 405798 319592
rect 200114 319472 200120 319524
rect 200172 319512 200178 319524
rect 303890 319512 303896 319524
rect 200172 319484 303896 319512
rect 200172 319472 200178 319484
rect 303890 319472 303896 319484
rect 303948 319472 303954 319524
rect 357710 319472 357716 319524
rect 357768 319512 357774 319524
rect 432046 319512 432052 319524
rect 357768 319484 432052 319512
rect 357768 319472 357774 319484
rect 432046 319472 432052 319484
rect 432104 319472 432110 319524
rect 84194 319404 84200 319456
rect 84252 319444 84258 319456
rect 276198 319444 276204 319456
rect 84252 319416 276204 319444
rect 84252 319404 84258 319416
rect 276198 319404 276204 319416
rect 276256 319404 276262 319456
rect 381446 319404 381452 319456
rect 381504 319444 381510 319456
rect 532694 319444 532700 319456
rect 381504 319416 532700 319444
rect 381504 319404 381510 319416
rect 532694 319404 532700 319416
rect 532752 319404 532758 319456
rect 197354 318180 197360 318232
rect 197412 318220 197418 318232
rect 302602 318220 302608 318232
rect 197412 318192 302608 318220
rect 197412 318180 197418 318192
rect 302602 318180 302608 318192
rect 302660 318180 302666 318232
rect 355042 318180 355048 318232
rect 355100 318220 355106 318232
rect 419534 318220 419540 318232
rect 355100 318192 419540 318220
rect 355100 318180 355106 318192
rect 419534 318180 419540 318192
rect 419592 318180 419598 318232
rect 184934 318112 184940 318164
rect 184992 318152 184998 318164
rect 299658 318152 299664 318164
rect 184992 318124 299664 318152
rect 184992 318112 184998 318124
rect 299658 318112 299664 318124
rect 299716 318112 299722 318164
rect 361850 318112 361856 318164
rect 361908 318152 361914 318164
rect 448606 318152 448612 318164
rect 361908 318124 448612 318152
rect 361908 318112 361914 318124
rect 448606 318112 448612 318124
rect 448664 318112 448670 318164
rect 93854 318044 93860 318096
rect 93912 318084 93918 318096
rect 279050 318084 279056 318096
rect 93912 318056 279056 318084
rect 93912 318044 93918 318056
rect 279050 318044 279056 318056
rect 279108 318044 279114 318096
rect 303614 318044 303620 318096
rect 303672 318084 303678 318096
rect 327442 318084 327448 318096
rect 303672 318056 327448 318084
rect 303672 318044 303678 318056
rect 327442 318044 327448 318056
rect 327500 318044 327506 318096
rect 382458 318044 382464 318096
rect 382516 318084 382522 318096
rect 539594 318084 539600 318096
rect 382516 318056 539600 318084
rect 382516 318044 382522 318056
rect 539594 318044 539600 318056
rect 539652 318044 539658 318096
rect 218054 316820 218060 316872
rect 218112 316860 218118 316872
rect 307938 316860 307944 316872
rect 218112 316832 307944 316860
rect 218112 316820 218118 316832
rect 307938 316820 307944 316832
rect 307996 316820 308002 316872
rect 349430 316820 349436 316872
rect 349488 316860 349494 316872
rect 398834 316860 398840 316872
rect 349488 316832 398840 316860
rect 349488 316820 349494 316832
rect 398834 316820 398840 316832
rect 398892 316820 398898 316872
rect 193214 316752 193220 316804
rect 193272 316792 193278 316804
rect 301130 316792 301136 316804
rect 193272 316764 301136 316792
rect 193272 316752 193278 316764
rect 301130 316752 301136 316764
rect 301188 316752 301194 316804
rect 356422 316752 356428 316804
rect 356480 316792 356486 316804
rect 423674 316792 423680 316804
rect 356480 316764 423680 316792
rect 356480 316752 356486 316764
rect 423674 316752 423680 316764
rect 423732 316752 423738 316804
rect 60734 316684 60740 316736
rect 60792 316724 60798 316736
rect 60792 316696 263594 316724
rect 60792 316684 60798 316696
rect 263566 316656 263594 316696
rect 263870 316684 263876 316736
rect 263928 316724 263934 316736
rect 264054 316724 264060 316736
rect 263928 316696 264060 316724
rect 263928 316684 263934 316696
rect 264054 316684 264060 316696
rect 264112 316684 264118 316736
rect 338666 316684 338672 316736
rect 338724 316724 338730 316736
rect 349246 316724 349252 316736
rect 338724 316696 349252 316724
rect 338724 316684 338730 316696
rect 349246 316684 349252 316696
rect 349304 316684 349310 316736
rect 385586 316684 385592 316736
rect 385644 316724 385650 316736
rect 550634 316724 550640 316736
rect 385644 316696 550640 316724
rect 385644 316684 385650 316696
rect 550634 316684 550640 316696
rect 550692 316684 550698 316736
rect 270770 316656 270776 316668
rect 263566 316628 270776 316656
rect 270770 316616 270776 316628
rect 270828 316616 270834 316668
rect 211154 315392 211160 315444
rect 211212 315432 211218 315444
rect 306558 315432 306564 315444
rect 211212 315404 306564 315432
rect 211212 315392 211218 315404
rect 306558 315392 306564 315404
rect 306616 315392 306622 315444
rect 360930 315392 360936 315444
rect 360988 315432 360994 315444
rect 430574 315432 430580 315444
rect 360988 315404 430580 315432
rect 360988 315392 360994 315404
rect 430574 315392 430580 315404
rect 430632 315392 430638 315444
rect 128354 315324 128360 315376
rect 128412 315364 128418 315376
rect 287238 315364 287244 315376
rect 128412 315336 287244 315364
rect 128412 315324 128418 315336
rect 287238 315324 287244 315336
rect 287296 315324 287302 315376
rect 365898 315324 365904 315376
rect 365956 315364 365962 315376
rect 466454 315364 466460 315376
rect 365956 315336 466460 315364
rect 365956 315324 365962 315336
rect 466454 315324 466460 315336
rect 466512 315324 466518 315376
rect 66254 315256 66260 315308
rect 66312 315296 66318 315308
rect 272058 315296 272064 315308
rect 66312 315268 272064 315296
rect 66312 315256 66318 315268
rect 272058 315256 272064 315268
rect 272116 315256 272122 315308
rect 386782 315256 386788 315308
rect 386840 315296 386846 315308
rect 554774 315296 554780 315308
rect 386840 315268 554780 315296
rect 386840 315256 386846 315268
rect 554774 315256 554780 315268
rect 554832 315256 554838 315308
rect 229094 314032 229100 314084
rect 229152 314072 229158 314084
rect 310790 314072 310796 314084
rect 229152 314044 310796 314072
rect 229152 314032 229158 314044
rect 310790 314032 310796 314044
rect 310848 314032 310854 314084
rect 195974 313964 195980 314016
rect 196032 314004 196038 314016
rect 302510 314004 302516 314016
rect 196032 313976 302516 314004
rect 196032 313964 196038 313976
rect 302510 313964 302516 313976
rect 302568 313964 302574 314016
rect 368750 313964 368756 314016
rect 368808 314004 368814 314016
rect 481634 314004 481640 314016
rect 368808 313976 481640 314004
rect 368808 313964 368814 313976
rect 481634 313964 481640 313976
rect 481692 313964 481698 314016
rect 57974 313896 57980 313948
rect 58032 313936 58038 313948
rect 270494 313936 270500 313948
rect 58032 313908 270500 313936
rect 58032 313896 58038 313908
rect 270494 313896 270500 313908
rect 270552 313896 270558 313948
rect 343818 313896 343824 313948
rect 343876 313936 343882 313948
rect 372706 313936 372712 313948
rect 343876 313908 372712 313936
rect 343876 313896 343882 313908
rect 372706 313896 372712 313908
rect 372764 313896 372770 313948
rect 386690 313896 386696 313948
rect 386748 313936 386754 313948
rect 557534 313936 557540 313948
rect 386748 313908 557540 313936
rect 386748 313896 386754 313908
rect 557534 313896 557540 313908
rect 557592 313896 557598 313948
rect 282178 313216 282184 313268
rect 282236 313256 282242 313268
rect 580166 313256 580172 313268
rect 282236 313228 580172 313256
rect 282236 313216 282242 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 223574 312672 223580 312724
rect 223632 312712 223638 312724
rect 309410 312712 309416 312724
rect 223632 312684 309416 312712
rect 223632 312672 223638 312684
rect 309410 312672 309416 312684
rect 309468 312672 309474 312724
rect 135254 312604 135260 312656
rect 135312 312644 135318 312656
rect 287790 312644 287796 312656
rect 135312 312616 287796 312644
rect 135312 312604 135318 312616
rect 287790 312604 287796 312616
rect 287848 312604 287854 312656
rect 44174 312536 44180 312588
rect 44232 312576 44238 312588
rect 266630 312576 266636 312588
rect 44232 312548 266636 312576
rect 44232 312536 44238 312548
rect 266630 312536 266636 312548
rect 266688 312536 266694 312588
rect 353386 312536 353392 312588
rect 353444 312576 353450 312588
rect 416774 312576 416780 312588
rect 353444 312548 416780 312576
rect 353444 312536 353450 312548
rect 416774 312536 416780 312548
rect 416832 312536 416838 312588
rect 236086 311244 236092 311296
rect 236144 311284 236150 311296
rect 312078 311284 312084 311296
rect 236144 311256 312084 311284
rect 236144 311244 236150 311256
rect 312078 311244 312084 311256
rect 312136 311244 312142 311296
rect 347958 311244 347964 311296
rect 348016 311284 348022 311296
rect 389174 311284 389180 311296
rect 348016 311256 389180 311284
rect 348016 311244 348022 311256
rect 389174 311244 389180 311256
rect 389232 311244 389238 311296
rect 202874 311176 202880 311228
rect 202932 311216 202938 311228
rect 303982 311216 303988 311228
rect 202932 311188 303988 311216
rect 202932 311176 202938 311188
rect 303982 311176 303988 311188
rect 304040 311176 304046 311228
rect 357618 311176 357624 311228
rect 357676 311216 357682 311228
rect 434714 311216 434720 311228
rect 357676 311188 434720 311216
rect 357676 311176 357682 311188
rect 434714 311176 434720 311188
rect 434772 311176 434778 311228
rect 4798 311108 4804 311160
rect 4856 311148 4862 311160
rect 256878 311148 256884 311160
rect 4856 311120 256884 311148
rect 4856 311108 4862 311120
rect 256878 311108 256884 311120
rect 256936 311108 256942 311160
rect 388162 311108 388168 311160
rect 388220 311148 388226 311160
rect 561674 311148 561680 311160
rect 388220 311120 561680 311148
rect 388220 311108 388226 311120
rect 561674 311108 561680 311120
rect 561732 311108 561738 311160
rect 209774 309884 209780 309936
rect 209832 309924 209838 309936
rect 305178 309924 305184 309936
rect 209832 309896 305184 309924
rect 209832 309884 209838 309896
rect 305178 309884 305184 309896
rect 305236 309884 305242 309936
rect 350718 309884 350724 309936
rect 350776 309924 350782 309936
rect 402974 309924 402980 309936
rect 350776 309896 402980 309924
rect 350776 309884 350782 309896
rect 402974 309884 402980 309896
rect 403032 309884 403038 309936
rect 147674 309816 147680 309868
rect 147732 309856 147738 309868
rect 291470 309856 291476 309868
rect 147732 309828 291476 309856
rect 147732 309816 147738 309828
rect 291470 309816 291476 309828
rect 291528 309816 291534 309868
rect 364610 309816 364616 309868
rect 364668 309856 364674 309868
rect 459554 309856 459560 309868
rect 364668 309828 459560 309856
rect 364668 309816 364674 309828
rect 459554 309816 459560 309828
rect 459612 309816 459618 309868
rect 77294 309748 77300 309800
rect 77352 309788 77358 309800
rect 273898 309788 273904 309800
rect 77352 309760 273904 309788
rect 77352 309748 77358 309760
rect 273898 309748 273904 309760
rect 273956 309748 273962 309800
rect 388070 309748 388076 309800
rect 388128 309788 388134 309800
rect 564434 309788 564440 309800
rect 388128 309760 564440 309788
rect 388128 309748 388134 309760
rect 564434 309748 564440 309760
rect 564492 309748 564498 309800
rect 227714 308524 227720 308576
rect 227772 308564 227778 308576
rect 309318 308564 309324 308576
rect 227772 308536 309324 308564
rect 227772 308524 227778 308536
rect 309318 308524 309324 308536
rect 309376 308524 309382 308576
rect 143534 308456 143540 308508
rect 143592 308496 143598 308508
rect 289906 308496 289912 308508
rect 143592 308468 289912 308496
rect 143592 308456 143598 308468
rect 289906 308456 289912 308468
rect 289964 308456 289970 308508
rect 352098 308456 352104 308508
rect 352156 308496 352162 308508
rect 409874 308496 409880 308508
rect 352156 308468 409880 308496
rect 352156 308456 352162 308468
rect 409874 308456 409880 308468
rect 409932 308456 409938 308508
rect 18598 308388 18604 308440
rect 18656 308428 18662 308440
rect 258166 308428 258172 308440
rect 18656 308400 258172 308428
rect 18656 308388 18662 308400
rect 258166 308388 258172 308400
rect 258224 308388 258230 308440
rect 389542 308388 389548 308440
rect 389600 308428 389606 308440
rect 567838 308428 567844 308440
rect 389600 308400 567844 308428
rect 389600 308388 389606 308400
rect 567838 308388 567844 308400
rect 567896 308388 567902 308440
rect 245654 307164 245660 307216
rect 245712 307204 245718 307216
rect 313458 307204 313464 307216
rect 245712 307176 313464 307204
rect 245712 307164 245718 307176
rect 313458 307164 313464 307176
rect 313516 307164 313522 307216
rect 179414 307096 179420 307148
rect 179472 307136 179478 307148
rect 298186 307136 298192 307148
rect 179472 307108 298192 307136
rect 179472 307096 179478 307108
rect 298186 307096 298192 307108
rect 298244 307096 298250 307148
rect 356330 307096 356336 307148
rect 356388 307136 356394 307148
rect 427814 307136 427820 307148
rect 356388 307108 427820 307136
rect 356388 307096 356394 307108
rect 427814 307096 427820 307108
rect 427872 307096 427878 307148
rect 75914 307028 75920 307080
rect 75972 307068 75978 307080
rect 274910 307068 274916 307080
rect 75972 307040 274916 307068
rect 75972 307028 75978 307040
rect 274910 307028 274916 307040
rect 274968 307028 274974 307080
rect 345290 307028 345296 307080
rect 345348 307068 345354 307080
rect 378226 307068 378232 307080
rect 345348 307040 378232 307068
rect 345348 307028 345354 307040
rect 378226 307028 378232 307040
rect 378284 307028 378290 307080
rect 390922 307028 390928 307080
rect 390980 307068 390986 307080
rect 575474 307068 575480 307080
rect 390980 307040 575480 307068
rect 390980 307028 390986 307040
rect 575474 307028 575480 307040
rect 575532 307028 575538 307080
rect 2774 306212 2780 306264
rect 2832 306252 2838 306264
rect 4890 306252 4896 306264
rect 2832 306224 4896 306252
rect 2832 306212 2838 306224
rect 4890 306212 4896 306224
rect 4948 306212 4954 306264
rect 247034 305736 247040 305788
rect 247092 305776 247098 305788
rect 314838 305776 314844 305788
rect 247092 305748 314844 305776
rect 247092 305736 247098 305748
rect 314838 305736 314844 305748
rect 314896 305736 314902 305788
rect 353570 305736 353576 305788
rect 353628 305776 353634 305788
rect 415394 305776 415400 305788
rect 353628 305748 415400 305776
rect 353628 305736 353634 305748
rect 415394 305736 415400 305748
rect 415452 305736 415458 305788
rect 139394 305668 139400 305720
rect 139452 305708 139458 305720
rect 288618 305708 288624 305720
rect 139452 305680 288624 305708
rect 139452 305668 139458 305680
rect 288618 305668 288624 305680
rect 288676 305668 288682 305720
rect 367278 305668 367284 305720
rect 367336 305708 367342 305720
rect 473354 305708 473360 305720
rect 367336 305680 473360 305708
rect 367336 305668 367342 305680
rect 473354 305668 473360 305680
rect 473412 305668 473418 305720
rect 40034 305600 40040 305652
rect 40092 305640 40098 305652
rect 264238 305640 264244 305652
rect 40092 305612 264244 305640
rect 40092 305600 40098 305612
rect 264238 305600 264244 305612
rect 264296 305600 264302 305652
rect 339678 305600 339684 305652
rect 339736 305640 339742 305652
rect 353386 305640 353392 305652
rect 339736 305612 353392 305640
rect 339736 305600 339742 305612
rect 353386 305600 353392 305612
rect 353444 305600 353450 305652
rect 378410 305600 378416 305652
rect 378468 305640 378474 305652
rect 521654 305640 521660 305652
rect 378468 305612 521660 305640
rect 378468 305600 378474 305612
rect 521654 305600 521660 305612
rect 521712 305600 521718 305652
rect 201586 304376 201592 304428
rect 201644 304416 201650 304428
rect 303798 304416 303804 304428
rect 201644 304388 303804 304416
rect 201644 304376 201650 304388
rect 303798 304376 303804 304388
rect 303856 304376 303862 304428
rect 143626 304308 143632 304360
rect 143684 304348 143690 304360
rect 289170 304348 289176 304360
rect 143684 304320 289176 304348
rect 143684 304308 143690 304320
rect 289170 304308 289176 304320
rect 289228 304308 289234 304360
rect 354674 304308 354680 304360
rect 354732 304348 354738 304360
rect 423766 304348 423772 304360
rect 354732 304320 423772 304348
rect 354732 304308 354738 304320
rect 423766 304308 423772 304320
rect 423824 304308 423830 304360
rect 88334 304240 88340 304292
rect 88392 304280 88398 304292
rect 277762 304280 277768 304292
rect 88392 304252 277768 304280
rect 88392 304240 88398 304252
rect 277762 304240 277768 304252
rect 277820 304240 277826 304292
rect 372982 304240 372988 304292
rect 373040 304280 373046 304292
rect 495434 304280 495440 304292
rect 373040 304252 495440 304280
rect 373040 304240 373046 304252
rect 495434 304240 495440 304252
rect 495492 304240 495498 304292
rect 219434 303016 219440 303068
rect 219492 303056 219498 303068
rect 307846 303056 307852 303068
rect 219492 303028 307852 303056
rect 219492 303016 219498 303028
rect 307846 303016 307852 303028
rect 307904 303016 307910 303068
rect 146294 302948 146300 303000
rect 146352 302988 146358 303000
rect 291378 302988 291384 303000
rect 146352 302960 291384 302988
rect 146352 302948 146358 302960
rect 291378 302948 291384 302960
rect 291436 302948 291442 303000
rect 357526 302948 357532 303000
rect 357584 302988 357590 303000
rect 433334 302988 433340 303000
rect 357584 302960 433340 302988
rect 357584 302948 357590 302960
rect 433334 302948 433340 302960
rect 433392 302948 433398 303000
rect 27614 302880 27620 302932
rect 27672 302920 27678 302932
rect 262398 302920 262404 302932
rect 27672 302892 262404 302920
rect 27672 302880 27678 302892
rect 262398 302880 262404 302892
rect 262456 302880 262462 302932
rect 377398 302880 377404 302932
rect 377456 302920 377462 302932
rect 509234 302920 509240 302932
rect 377456 302892 509240 302920
rect 377456 302880 377462 302892
rect 509234 302880 509240 302892
rect 509292 302880 509298 302932
rect 230474 301588 230480 301640
rect 230532 301628 230538 301640
rect 310698 301628 310704 301640
rect 230532 301600 310704 301628
rect 230532 301588 230538 301600
rect 310698 301588 310704 301600
rect 310756 301588 310762 301640
rect 150434 301520 150440 301572
rect 150492 301560 150498 301572
rect 291286 301560 291292 301572
rect 150492 301532 291292 301560
rect 150492 301520 150498 301532
rect 291286 301520 291292 301532
rect 291344 301520 291350 301572
rect 358998 301520 359004 301572
rect 359056 301560 359062 301572
rect 437474 301560 437480 301572
rect 359056 301532 437480 301560
rect 359056 301520 359062 301532
rect 437474 301520 437480 301532
rect 437532 301520 437538 301572
rect 22738 301452 22744 301504
rect 22796 301492 22802 301504
rect 259730 301492 259736 301504
rect 22796 301464 259736 301492
rect 22796 301452 22802 301464
rect 259730 301452 259736 301464
rect 259788 301452 259794 301504
rect 378318 301452 378324 301504
rect 378376 301492 378382 301504
rect 520274 301492 520280 301504
rect 378376 301464 520280 301492
rect 378376 301452 378382 301464
rect 520274 301452 520280 301464
rect 520332 301452 520338 301504
rect 153194 300160 153200 300212
rect 153252 300200 153258 300212
rect 292758 300200 292764 300212
rect 153252 300172 292764 300200
rect 153252 300160 153258 300172
rect 292758 300160 292764 300172
rect 292816 300160 292822 300212
rect 358906 300160 358912 300212
rect 358964 300200 358970 300212
rect 440326 300200 440332 300212
rect 358964 300172 440332 300200
rect 358964 300160 358970 300172
rect 440326 300160 440332 300172
rect 440384 300160 440390 300212
rect 110506 300092 110512 300144
rect 110564 300132 110570 300144
rect 283282 300132 283288 300144
rect 110564 300104 283288 300132
rect 110564 300092 110570 300104
rect 283282 300092 283288 300104
rect 283340 300092 283346 300144
rect 381170 300092 381176 300144
rect 381228 300132 381234 300144
rect 531314 300132 531320 300144
rect 381228 300104 531320 300132
rect 381228 300092 381234 300104
rect 531314 300092 531320 300104
rect 531372 300092 531378 300144
rect 567930 299412 567936 299464
rect 567988 299452 567994 299464
rect 579614 299452 579620 299464
rect 567988 299424 579620 299452
rect 567988 299412 567994 299424
rect 579614 299412 579620 299424
rect 579672 299412 579678 299464
rect 157334 298800 157340 298852
rect 157392 298840 157398 298852
rect 292666 298840 292672 298852
rect 157392 298812 292672 298840
rect 157392 298800 157398 298812
rect 292666 298800 292672 298812
rect 292724 298800 292730 298852
rect 360378 298800 360384 298852
rect 360436 298840 360442 298852
rect 444374 298840 444380 298852
rect 360436 298812 444380 298840
rect 360436 298800 360442 298812
rect 444374 298800 444380 298812
rect 444432 298800 444438 298852
rect 26234 298732 26240 298784
rect 26292 298772 26298 298784
rect 261478 298772 261484 298784
rect 26292 298744 261484 298772
rect 26292 298732 26298 298744
rect 261478 298732 261484 298744
rect 261536 298732 261542 298784
rect 385034 298732 385040 298784
rect 385092 298772 385098 298784
rect 552014 298772 552020 298784
rect 385092 298744 552020 298772
rect 385092 298732 385098 298744
rect 552014 298732 552020 298744
rect 552072 298732 552078 298784
rect 255314 297508 255320 297560
rect 255372 297548 255378 297560
rect 316218 297548 316224 297560
rect 255372 297520 316224 297548
rect 255372 297508 255378 297520
rect 316218 297508 316224 297520
rect 316276 297508 316282 297560
rect 126974 297440 126980 297492
rect 127032 297480 127038 297492
rect 285950 297480 285956 297492
rect 127032 297452 285956 297480
rect 127032 297440 127038 297452
rect 285950 297440 285956 297452
rect 286008 297440 286014 297492
rect 361666 297440 361672 297492
rect 361724 297480 361730 297492
rect 451274 297480 451280 297492
rect 361724 297452 451280 297480
rect 361724 297440 361730 297452
rect 451274 297440 451280 297452
rect 451332 297440 451338 297492
rect 102134 297372 102140 297424
rect 102192 297412 102198 297424
rect 280338 297412 280344 297424
rect 102192 297384 280344 297412
rect 102192 297372 102198 297384
rect 280338 297372 280344 297384
rect 280396 297372 280402 297424
rect 390646 297372 390652 297424
rect 390704 297412 390710 297424
rect 572070 297412 572076 297424
rect 390704 297384 572076 297412
rect 390704 297372 390710 297384
rect 572070 297372 572076 297384
rect 572128 297372 572134 297424
rect 165614 296012 165620 296064
rect 165672 296052 165678 296064
rect 295426 296052 295432 296064
rect 165672 296024 295432 296052
rect 165672 296012 165678 296024
rect 295426 296012 295432 296024
rect 295484 296012 295490 296064
rect 363230 296012 363236 296064
rect 363288 296052 363294 296064
rect 455414 296052 455420 296064
rect 363288 296024 455420 296052
rect 363288 296012 363294 296024
rect 455414 296012 455420 296024
rect 455472 296012 455478 296064
rect 35894 295944 35900 295996
rect 35952 295984 35958 295996
rect 265250 295984 265256 295996
rect 35952 295956 265256 295984
rect 35952 295944 35958 295956
rect 265250 295944 265256 295956
rect 265308 295944 265314 295996
rect 365806 295944 365812 295996
rect 365864 295984 365870 295996
rect 470594 295984 470600 295996
rect 365864 295956 470600 295984
rect 365864 295944 365870 295956
rect 470594 295944 470600 295956
rect 470652 295944 470658 295996
rect 176654 294652 176660 294704
rect 176712 294692 176718 294704
rect 297450 294692 297456 294704
rect 176712 294664 297456 294692
rect 176712 294652 176718 294664
rect 297450 294652 297456 294664
rect 297508 294652 297514 294704
rect 363138 294652 363144 294704
rect 363196 294692 363202 294704
rect 458174 294692 458180 294704
rect 363196 294664 458180 294692
rect 363196 294652 363202 294664
rect 458174 294652 458180 294664
rect 458232 294652 458238 294704
rect 20714 294584 20720 294636
rect 20772 294624 20778 294636
rect 261110 294624 261116 294636
rect 20772 294596 261116 294624
rect 20772 294584 20778 294596
rect 261110 294584 261116 294596
rect 261168 294584 261174 294636
rect 296714 294584 296720 294636
rect 296772 294624 296778 294636
rect 325878 294624 325884 294636
rect 296772 294596 325884 294624
rect 296772 294584 296778 294596
rect 325878 294584 325884 294596
rect 325936 294584 325942 294636
rect 371234 294584 371240 294636
rect 371292 294624 371298 294636
rect 490006 294624 490012 294636
rect 371292 294596 490012 294624
rect 371292 294584 371298 294596
rect 490006 294584 490012 294596
rect 490064 294584 490070 294636
rect 3050 293904 3056 293956
rect 3108 293944 3114 293956
rect 221458 293944 221464 293956
rect 3108 293916 221464 293944
rect 3108 293904 3114 293916
rect 221458 293904 221464 293916
rect 221516 293904 221522 293956
rect 369118 293292 369124 293344
rect 369176 293332 369182 293344
rect 465166 293332 465172 293344
rect 369176 293304 465172 293332
rect 369176 293292 369182 293304
rect 465166 293292 465172 293304
rect 465224 293292 465230 293344
rect 215294 293224 215300 293276
rect 215352 293264 215358 293276
rect 306466 293264 306472 293276
rect 215352 293236 306472 293264
rect 215352 293224 215358 293236
rect 306466 293224 306472 293236
rect 306524 293224 306530 293276
rect 375466 293224 375472 293276
rect 375524 293264 375530 293276
rect 506474 293264 506480 293276
rect 375524 293236 506480 293264
rect 375524 293224 375530 293236
rect 506474 293224 506480 293236
rect 506532 293224 506538 293276
rect 299658 292000 299664 292052
rect 299716 292040 299722 292052
rect 327350 292040 327356 292052
rect 299716 292012 327356 292040
rect 299716 292000 299722 292012
rect 327350 292000 327356 292012
rect 327408 292000 327414 292052
rect 183554 291864 183560 291916
rect 183612 291904 183618 291916
rect 299566 291904 299572 291916
rect 183612 291876 299572 291904
rect 183612 291864 183618 291876
rect 299566 291864 299572 291876
rect 299624 291864 299630 291916
rect 367462 291864 367468 291916
rect 367520 291904 367526 291916
rect 476114 291904 476120 291916
rect 367520 291876 476120 291904
rect 367520 291864 367526 291876
rect 476114 291864 476120 291876
rect 476172 291864 476178 291916
rect 28994 291796 29000 291848
rect 29052 291836 29058 291848
rect 263870 291836 263876 291848
rect 29052 291808 263876 291836
rect 29052 291796 29058 291808
rect 263870 291796 263876 291808
rect 263928 291796 263934 291848
rect 342530 291796 342536 291848
rect 342588 291836 342594 291848
rect 367278 291836 367284 291848
rect 342588 291808 367284 291836
rect 342588 291796 342594 291808
rect 367278 291796 367284 291808
rect 367336 291796 367342 291848
rect 379606 291796 379612 291848
rect 379664 291836 379670 291848
rect 524414 291836 524420 291848
rect 379664 291808 524420 291836
rect 379664 291796 379670 291808
rect 524414 291796 524420 291808
rect 524472 291796 524478 291848
rect 190454 290504 190460 290556
rect 190512 290544 190518 290556
rect 301038 290544 301044 290556
rect 190512 290516 301044 290544
rect 190512 290504 190518 290516
rect 301038 290504 301044 290516
rect 301096 290504 301102 290556
rect 370038 290504 370044 290556
rect 370096 290544 370102 290556
rect 484394 290544 484400 290556
rect 370096 290516 484400 290544
rect 370096 290504 370102 290516
rect 484394 290504 484400 290516
rect 484452 290504 484458 290556
rect 114554 290436 114560 290488
rect 114612 290476 114618 290488
rect 283190 290476 283196 290488
rect 114612 290448 283196 290476
rect 114612 290436 114618 290448
rect 283190 290436 283196 290448
rect 283248 290436 283254 290488
rect 383746 290436 383752 290488
rect 383804 290476 383810 290488
rect 542354 290476 542360 290488
rect 383804 290448 542360 290476
rect 383804 290436 383810 290448
rect 542354 290436 542360 290448
rect 542412 290436 542418 290488
rect 193306 289144 193312 289196
rect 193364 289184 193370 289196
rect 302418 289184 302424 289196
rect 193364 289156 302424 289184
rect 193364 289144 193370 289156
rect 302418 289144 302424 289156
rect 302476 289144 302482 289196
rect 16574 289076 16580 289128
rect 16632 289116 16638 289128
rect 256142 289116 256148 289128
rect 16632 289088 256148 289116
rect 16632 289076 16638 289088
rect 256142 289076 256148 289088
rect 256200 289076 256206 289128
rect 369946 289076 369952 289128
rect 370004 289116 370010 289128
rect 488534 289116 488540 289128
rect 370004 289088 488540 289116
rect 370004 289076 370010 289088
rect 488534 289076 488540 289088
rect 488592 289076 488598 289128
rect 129734 287716 129740 287768
rect 129792 287756 129798 287768
rect 287146 287756 287152 287768
rect 129792 287728 287152 287756
rect 129792 287716 129798 287728
rect 287146 287716 287152 287728
rect 287204 287716 287210 287768
rect 60826 287648 60832 287700
rect 60884 287688 60890 287700
rect 269758 287688 269764 287700
rect 60884 287660 269764 287688
rect 60884 287648 60890 287660
rect 269758 287648 269764 287660
rect 269816 287648 269822 287700
rect 345658 287648 345664 287700
rect 345716 287688 345722 287700
rect 371234 287688 371240 287700
rect 345716 287660 371240 287688
rect 345716 287648 345722 287660
rect 371234 287648 371240 287660
rect 371292 287648 371298 287700
rect 371418 287648 371424 287700
rect 371476 287688 371482 287700
rect 491294 287688 491300 287700
rect 371476 287660 491300 287688
rect 371476 287648 371482 287660
rect 491294 287648 491300 287660
rect 491352 287648 491358 287700
rect 208394 286356 208400 286408
rect 208452 286396 208458 286408
rect 305086 286396 305092 286408
rect 208452 286368 305092 286396
rect 208452 286356 208458 286368
rect 305086 286356 305092 286368
rect 305144 286356 305150 286408
rect 96614 286288 96620 286340
rect 96672 286328 96678 286340
rect 278958 286328 278964 286340
rect 96672 286300 278964 286328
rect 96672 286288 96678 286300
rect 278958 286288 278964 286300
rect 279016 286288 279022 286340
rect 372890 286288 372896 286340
rect 372948 286328 372954 286340
rect 498286 286328 498292 286340
rect 372948 286300 498292 286328
rect 372948 286288 372954 286300
rect 498286 286288 498292 286300
rect 498344 286288 498350 286340
rect 307754 285132 307760 285184
rect 307812 285172 307818 285184
rect 328822 285172 328828 285184
rect 307812 285144 328828 285172
rect 307812 285132 307818 285144
rect 328822 285132 328828 285144
rect 328880 285132 328886 285184
rect 222194 284996 222200 285048
rect 222252 285036 222258 285048
rect 308030 285036 308036 285048
rect 222252 285008 308036 285036
rect 222252 284996 222258 285008
rect 308030 284996 308036 285008
rect 308088 284996 308094 285048
rect 78674 284928 78680 284980
rect 78732 284968 78738 284980
rect 274818 284968 274824 284980
rect 78732 284940 274824 284968
rect 78732 284928 78738 284940
rect 274818 284928 274824 284940
rect 274876 284928 274882 284980
rect 343726 284928 343732 284980
rect 343784 284968 343790 284980
rect 374086 284968 374092 284980
rect 343784 284940 374092 284968
rect 343784 284928 343790 284940
rect 374086 284928 374092 284940
rect 374144 284928 374150 284980
rect 374362 284928 374368 284980
rect 374420 284968 374426 284980
rect 502334 284968 502340 284980
rect 374420 284940 502340 284968
rect 374420 284928 374426 284940
rect 502334 284928 502340 284940
rect 502392 284928 502398 284980
rect 226334 283636 226340 283688
rect 226392 283676 226398 283688
rect 309226 283676 309232 283688
rect 226392 283648 309232 283676
rect 226392 283636 226398 283648
rect 309226 283636 309232 283648
rect 309284 283636 309290 283688
rect 89714 283568 89720 283620
rect 89772 283608 89778 283620
rect 277670 283608 277676 283620
rect 89772 283580 277676 283608
rect 89772 283568 89778 283580
rect 277670 283568 277676 283580
rect 277728 283568 277734 283620
rect 374270 283568 374276 283620
rect 374328 283608 374334 283620
rect 506566 283608 506572 283620
rect 374328 283580 506572 283608
rect 374328 283568 374334 283580
rect 506566 283568 506572 283580
rect 506624 283568 506630 283620
rect 133874 282140 133880 282192
rect 133932 282180 133938 282192
rect 287330 282180 287336 282192
rect 133932 282152 287336 282180
rect 133932 282140 133938 282152
rect 287330 282140 287336 282152
rect 287388 282140 287394 282192
rect 376938 282140 376944 282192
rect 376996 282180 377002 282192
rect 516134 282180 516140 282192
rect 376996 282152 516140 282180
rect 376996 282140 377002 282152
rect 516134 282140 516140 282152
rect 516192 282140 516198 282192
rect 233234 280848 233240 280900
rect 233292 280888 233298 280900
rect 310606 280888 310612 280900
rect 233292 280860 310612 280888
rect 233292 280848 233298 280860
rect 310606 280848 310612 280860
rect 310664 280848 310670 280900
rect 64874 280780 64880 280832
rect 64932 280820 64938 280832
rect 268378 280820 268384 280832
rect 64932 280792 268384 280820
rect 64932 280780 64938 280792
rect 268378 280780 268384 280792
rect 268436 280780 268442 280832
rect 381078 280780 381084 280832
rect 381136 280820 381142 280832
rect 534074 280820 534080 280832
rect 381136 280792 534080 280820
rect 381136 280780 381142 280792
rect 534074 280780 534080 280792
rect 534132 280780 534138 280832
rect 240134 279488 240140 279540
rect 240192 279528 240198 279540
rect 311986 279528 311992 279540
rect 240192 279500 311992 279528
rect 240192 279488 240198 279500
rect 311986 279488 311992 279500
rect 312044 279488 312050 279540
rect 8938 279420 8944 279472
rect 8996 279460 9002 279472
rect 256786 279460 256792 279472
rect 8996 279432 256792 279460
rect 8996 279420 9002 279432
rect 256786 279420 256792 279432
rect 256844 279420 256850 279472
rect 346670 279420 346676 279472
rect 346728 279460 346734 279472
rect 382458 279460 382464 279472
rect 346728 279432 382464 279460
rect 346728 279420 346734 279432
rect 382458 279420 382464 279432
rect 382516 279420 382522 279472
rect 382550 279420 382556 279472
rect 382608 279460 382614 279472
rect 538214 279460 538220 279472
rect 382608 279432 538220 279460
rect 382608 279420 382614 279432
rect 538214 279420 538220 279432
rect 538272 279420 538278 279472
rect 314654 278196 314660 278248
rect 314712 278236 314718 278248
rect 330018 278236 330024 278248
rect 314712 278208 330024 278236
rect 314712 278196 314718 278208
rect 330018 278196 330024 278208
rect 330076 278196 330082 278248
rect 251174 278060 251180 278112
rect 251232 278100 251238 278112
rect 315022 278100 315028 278112
rect 251232 278072 315028 278100
rect 251232 278060 251238 278072
rect 315022 278060 315028 278072
rect 315080 278060 315086 278112
rect 7558 277992 7564 278044
rect 7616 278032 7622 278044
rect 256970 278032 256976 278044
rect 7616 278004 256976 278032
rect 7616 277992 7622 278004
rect 256970 277992 256976 278004
rect 257028 277992 257034 278044
rect 346578 277992 346584 278044
rect 346636 278032 346642 278044
rect 385034 278032 385040 278044
rect 346636 278004 385040 278032
rect 346636 277992 346642 278004
rect 385034 277992 385040 278004
rect 385092 277992 385098 278044
rect 385310 277992 385316 278044
rect 385368 278032 385374 278044
rect 547966 278032 547972 278044
rect 385368 278004 547972 278032
rect 385368 277992 385374 278004
rect 547966 277992 547972 278004
rect 548024 277992 548030 278044
rect 151814 276632 151820 276684
rect 151872 276672 151878 276684
rect 291562 276672 291568 276684
rect 151872 276644 291568 276672
rect 151872 276632 151878 276644
rect 291562 276632 291568 276644
rect 291620 276632 291626 276684
rect 386598 276632 386604 276684
rect 386656 276672 386662 276684
rect 556154 276672 556160 276684
rect 386656 276644 556160 276672
rect 386656 276632 386662 276644
rect 556154 276632 556160 276644
rect 556212 276632 556218 276684
rect 162854 275340 162860 275392
rect 162912 275380 162918 275392
rect 294138 275380 294144 275392
rect 162912 275352 294144 275380
rect 162912 275340 162918 275352
rect 294138 275340 294144 275352
rect 294196 275340 294202 275392
rect 81434 275272 81440 275324
rect 81492 275312 81498 275324
rect 276106 275312 276112 275324
rect 81492 275284 276112 275312
rect 81492 275272 81498 275284
rect 276106 275272 276112 275284
rect 276164 275272 276170 275324
rect 387978 275272 387984 275324
rect 388036 275312 388042 275324
rect 563054 275312 563060 275324
rect 388036 275284 563060 275312
rect 388036 275272 388042 275284
rect 563054 275272 563060 275284
rect 563112 275272 563118 275324
rect 166994 273980 167000 274032
rect 167052 274020 167058 274032
rect 295610 274020 295616 274032
rect 167052 273992 295616 274020
rect 167052 273980 167058 273992
rect 295610 273980 295616 273992
rect 295668 273980 295674 274032
rect 99374 273912 99380 273964
rect 99432 273952 99438 273964
rect 280246 273952 280252 273964
rect 99432 273924 280252 273952
rect 99432 273912 99438 273924
rect 280246 273912 280252 273924
rect 280304 273912 280310 273964
rect 389450 273912 389456 273964
rect 389508 273952 389514 273964
rect 569954 273952 569960 273964
rect 389508 273924 569960 273952
rect 389508 273912 389514 273924
rect 569954 273912 569960 273924
rect 570012 273912 570018 273964
rect 431218 273164 431224 273216
rect 431276 273204 431282 273216
rect 579890 273204 579896 273216
rect 431276 273176 579896 273204
rect 431276 273164 431282 273176
rect 579890 273164 579896 273176
rect 579948 273164 579954 273216
rect 169754 272552 169760 272604
rect 169812 272592 169818 272604
rect 296898 272592 296904 272604
rect 169812 272564 296904 272592
rect 169812 272552 169818 272564
rect 296898 272552 296904 272564
rect 296956 272552 296962 272604
rect 106274 272484 106280 272536
rect 106332 272524 106338 272536
rect 281810 272524 281816 272536
rect 106332 272496 281816 272524
rect 106332 272484 106338 272496
rect 281810 272484 281816 272496
rect 281868 272484 281874 272536
rect 353478 272484 353484 272536
rect 353536 272524 353542 272536
rect 414014 272524 414020 272536
rect 353536 272496 414020 272524
rect 353536 272484 353542 272496
rect 414014 272484 414020 272496
rect 414072 272484 414078 272536
rect 173894 271124 173900 271176
rect 173952 271164 173958 271176
rect 296806 271164 296812 271176
rect 173952 271136 296812 271164
rect 173952 271124 173958 271136
rect 296806 271124 296812 271136
rect 296864 271124 296870 271176
rect 347866 271124 347872 271176
rect 347924 271164 347930 271176
rect 390646 271164 390652 271176
rect 347924 271136 390652 271164
rect 347924 271124 347930 271136
rect 390646 271124 390652 271136
rect 390704 271124 390710 271176
rect 390830 271124 390836 271176
rect 390888 271164 390894 271176
rect 574738 271164 574744 271176
rect 390888 271136 574744 271164
rect 390888 271124 390894 271136
rect 574738 271124 574744 271136
rect 574796 271124 574802 271176
rect 180794 269832 180800 269884
rect 180852 269872 180858 269884
rect 298278 269872 298284 269884
rect 180852 269844 298284 269872
rect 180852 269832 180858 269844
rect 298278 269832 298284 269844
rect 298336 269832 298342 269884
rect 354950 269832 354956 269884
rect 355008 269872 355014 269884
rect 420914 269872 420920 269884
rect 355008 269844 420920 269872
rect 355008 269832 355014 269844
rect 420914 269832 420920 269844
rect 420972 269832 420978 269884
rect 63494 269764 63500 269816
rect 63552 269804 63558 269816
rect 271966 269804 271972 269816
rect 63552 269776 271972 269804
rect 63552 269764 63558 269776
rect 271966 269764 271972 269776
rect 272024 269764 272030 269816
rect 341518 269764 341524 269816
rect 341576 269804 341582 269816
rect 354674 269804 354680 269816
rect 341576 269776 354680 269804
rect 341576 269764 341582 269776
rect 354674 269764 354680 269776
rect 354732 269764 354738 269816
rect 385218 269764 385224 269816
rect 385276 269804 385282 269816
rect 549254 269804 549260 269816
rect 385276 269776 549260 269804
rect 385276 269764 385282 269776
rect 549254 269764 549260 269776
rect 549312 269764 549318 269816
rect 185026 268404 185032 268456
rect 185084 268444 185090 268456
rect 298738 268444 298744 268456
rect 185084 268416 298744 268444
rect 185084 268404 185090 268416
rect 298738 268404 298744 268416
rect 298796 268404 298802 268456
rect 70394 268336 70400 268388
rect 70452 268376 70458 268388
rect 273530 268376 273536 268388
rect 70452 268348 273536 268376
rect 70452 268336 70458 268348
rect 273530 268336 273536 268348
rect 273588 268336 273594 268388
rect 360286 268336 360292 268388
rect 360344 268376 360350 268388
rect 445754 268376 445760 268388
rect 360344 268348 445760 268376
rect 360344 268336 360350 268348
rect 445754 268336 445760 268348
rect 445812 268336 445818 268388
rect 3510 267656 3516 267708
rect 3568 267696 3574 267708
rect 232498 267696 232504 267708
rect 3568 267668 232504 267696
rect 3568 267656 3574 267668
rect 232498 267656 232504 267668
rect 232556 267656 232562 267708
rect 234706 266976 234712 267028
rect 234764 267016 234770 267028
rect 310882 267016 310888 267028
rect 234764 266988 310888 267016
rect 234764 266976 234770 266988
rect 310882 266976 310888 266988
rect 310940 266976 310946 267028
rect 361574 266976 361580 267028
rect 361632 267016 361638 267028
rect 452654 267016 452660 267028
rect 361632 266988 452660 267016
rect 361632 266976 361638 266988
rect 452654 266976 452660 266988
rect 452712 266976 452718 267028
rect 187694 265616 187700 265668
rect 187752 265656 187758 265668
rect 300946 265656 300952 265668
rect 187752 265628 300952 265656
rect 187752 265616 187758 265628
rect 300946 265616 300952 265628
rect 301004 265616 301010 265668
rect 363046 265616 363052 265668
rect 363104 265656 363110 265668
rect 456886 265656 456892 265668
rect 363104 265628 456892 265656
rect 363104 265616 363110 265628
rect 456886 265616 456892 265628
rect 456944 265616 456950 265668
rect 191834 264188 191840 264240
rect 191892 264228 191898 264240
rect 301222 264228 301228 264240
rect 191892 264200 301228 264228
rect 191892 264188 191898 264200
rect 301222 264188 301228 264200
rect 301280 264188 301286 264240
rect 364518 264188 364524 264240
rect 364576 264228 364582 264240
rect 463694 264228 463700 264240
rect 364576 264200 463700 264228
rect 364576 264188 364582 264200
rect 463694 264188 463700 264200
rect 463752 264188 463758 264240
rect 198734 262896 198740 262948
rect 198792 262936 198798 262948
rect 302326 262936 302332 262948
rect 198792 262908 302332 262936
rect 198792 262896 198798 262908
rect 302326 262896 302332 262908
rect 302384 262896 302390 262948
rect 41414 262828 41420 262880
rect 41472 262868 41478 262880
rect 266538 262868 266544 262880
rect 41472 262840 266544 262868
rect 41472 262828 41478 262840
rect 266538 262828 266544 262840
rect 266596 262828 266602 262880
rect 367370 262828 367376 262880
rect 367428 262868 367434 262880
rect 473446 262868 473452 262880
rect 367428 262840 473452 262868
rect 367428 262828 367434 262840
rect 473446 262828 473452 262840
rect 473504 262828 473510 262880
rect 135346 261468 135352 261520
rect 135404 261508 135410 261520
rect 288526 261508 288532 261520
rect 135404 261480 288532 261508
rect 135404 261468 135410 261480
rect 288526 261468 288532 261480
rect 288584 261468 288590 261520
rect 368658 261468 368664 261520
rect 368716 261508 368722 261520
rect 477494 261508 477500 261520
rect 368716 261480 477500 261508
rect 368716 261468 368722 261480
rect 477494 261468 477500 261480
rect 477552 261468 477558 261520
rect 241514 260176 241520 260228
rect 241572 260216 241578 260228
rect 313366 260216 313372 260228
rect 241572 260188 313372 260216
rect 241572 260176 241578 260188
rect 313366 260176 313372 260188
rect 313424 260176 313430 260228
rect 52454 260108 52460 260160
rect 52512 260148 52518 260160
rect 269390 260148 269396 260160
rect 52512 260120 269396 260148
rect 52512 260108 52518 260120
rect 269390 260108 269396 260120
rect 269448 260108 269454 260160
rect 369854 260108 369860 260160
rect 369912 260148 369918 260160
rect 485774 260148 485780 260160
rect 369912 260120 485780 260148
rect 369912 260108 369918 260120
rect 485774 260108 485780 260120
rect 485832 260108 485838 260160
rect 407850 259360 407856 259412
rect 407908 259400 407914 259412
rect 579798 259400 579804 259412
rect 407908 259372 579804 259400
rect 407908 259360 407914 259372
rect 579798 259360 579804 259372
rect 579856 259360 579862 259412
rect 138014 258680 138020 258732
rect 138072 258720 138078 258732
rect 288710 258720 288716 258732
rect 138072 258692 288716 258720
rect 138072 258680 138078 258692
rect 288710 258680 288716 258692
rect 288768 258680 288774 258732
rect 354858 258680 354864 258732
rect 354916 258720 354922 258732
rect 418154 258720 418160 258732
rect 354916 258692 418160 258720
rect 354916 258680 354922 258692
rect 418154 258680 418160 258692
rect 418212 258680 418218 258732
rect 144914 257320 144920 257372
rect 144972 257360 144978 257372
rect 290090 257360 290096 257372
rect 144972 257332 290096 257360
rect 144972 257320 144978 257332
rect 290090 257320 290096 257332
rect 290148 257320 290154 257372
rect 371326 257320 371332 257372
rect 371384 257360 371390 257372
rect 492674 257360 492680 257372
rect 371384 257332 492680 257360
rect 371384 257320 371390 257332
rect 492674 257320 492680 257332
rect 492732 257320 492738 257372
rect 151906 255960 151912 256012
rect 151964 256000 151970 256012
rect 292942 256000 292948 256012
rect 151964 255972 292948 256000
rect 151964 255960 151970 255972
rect 292942 255960 292948 255972
rect 293000 255960 293006 256012
rect 372798 255960 372804 256012
rect 372856 256000 372862 256012
rect 499574 256000 499580 256012
rect 372856 255972 499580 256000
rect 372856 255960 372862 255972
rect 499574 255960 499580 255972
rect 499632 255960 499638 256012
rect 3142 255212 3148 255264
rect 3200 255252 3206 255264
rect 14550 255252 14556 255264
rect 3200 255224 14556 255252
rect 3200 255212 3206 255224
rect 14550 255212 14556 255224
rect 14608 255212 14614 255264
rect 69014 254532 69020 254584
rect 69072 254572 69078 254584
rect 271230 254572 271236 254584
rect 69072 254544 271236 254572
rect 69072 254532 69078 254544
rect 271230 254532 271236 254544
rect 271288 254532 271294 254584
rect 374178 254532 374184 254584
rect 374236 254572 374242 254584
rect 503714 254572 503720 254584
rect 374236 254544 503720 254572
rect 374236 254532 374242 254544
rect 503714 254532 503720 254544
rect 503772 254532 503778 254584
rect 82814 253172 82820 253224
rect 82872 253212 82878 253224
rect 275278 253212 275284 253224
rect 82872 253184 275284 253212
rect 82872 253172 82878 253184
rect 275278 253172 275284 253184
rect 275336 253172 275342 253224
rect 375374 253172 375380 253224
rect 375432 253212 375438 253224
rect 510614 253212 510620 253224
rect 375432 253184 510620 253212
rect 375432 253172 375438 253184
rect 510614 253172 510620 253184
rect 510672 253172 510678 253224
rect 100754 251812 100760 251864
rect 100812 251852 100818 251864
rect 279418 251852 279424 251864
rect 100812 251824 279424 251852
rect 100812 251812 100818 251824
rect 279418 251812 279424 251824
rect 279476 251812 279482 251864
rect 376846 251812 376852 251864
rect 376904 251852 376910 251864
rect 517514 251852 517520 251864
rect 376904 251824 517520 251852
rect 376904 251812 376910 251824
rect 517514 251812 517520 251824
rect 517572 251812 517578 251864
rect 118694 250452 118700 250504
rect 118752 250492 118758 250504
rect 284570 250492 284576 250504
rect 118752 250464 284576 250492
rect 118752 250452 118758 250464
rect 284570 250452 284576 250464
rect 284628 250452 284634 250504
rect 379514 250452 379520 250504
rect 379572 250492 379578 250504
rect 528554 250492 528560 250504
rect 379572 250464 528560 250492
rect 379572 250452 379578 250464
rect 528554 250452 528560 250464
rect 528612 250452 528618 250504
rect 2774 249024 2780 249076
rect 2832 249064 2838 249076
rect 256050 249064 256056 249076
rect 2832 249036 256056 249064
rect 2832 249024 2838 249036
rect 256050 249024 256056 249036
rect 256108 249024 256114 249076
rect 380986 249024 380992 249076
rect 381044 249064 381050 249076
rect 535454 249064 535460 249076
rect 381044 249036 535460 249064
rect 381044 249024 381050 249036
rect 535454 249024 535460 249036
rect 535512 249024 535518 249076
rect 48314 247664 48320 247716
rect 48372 247704 48378 247716
rect 267918 247704 267924 247716
rect 48372 247676 267924 247704
rect 48372 247664 48378 247676
rect 267918 247664 267924 247676
rect 267976 247664 267982 247716
rect 383654 247664 383660 247716
rect 383712 247704 383718 247716
rect 546494 247704 546500 247716
rect 383712 247676 546500 247704
rect 383712 247664 383718 247676
rect 546494 247664 546500 247676
rect 546552 247664 546558 247716
rect 59354 246304 59360 246356
rect 59412 246344 59418 246356
rect 270586 246344 270592 246356
rect 59412 246316 270592 246344
rect 59412 246304 59418 246316
rect 270586 246304 270592 246316
rect 270644 246304 270650 246356
rect 385126 246304 385132 246356
rect 385184 246344 385190 246356
rect 553394 246344 553400 246356
rect 385184 246316 553400 246344
rect 385184 246304 385190 246316
rect 553394 246304 553400 246316
rect 553452 246304 553458 246356
rect 422938 245556 422944 245608
rect 422996 245596 423002 245608
rect 580166 245596 580172 245608
rect 422996 245568 580172 245596
rect 422996 245556 423002 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 62114 244876 62120 244928
rect 62172 244916 62178 244928
rect 270862 244916 270868 244928
rect 62172 244888 270868 244916
rect 62172 244876 62178 244888
rect 270862 244876 270868 244888
rect 270920 244876 270926 244928
rect 354766 244876 354772 244928
rect 354824 244916 354830 244928
rect 422294 244916 422300 244928
rect 354824 244888 422300 244916
rect 354824 244876 354830 244888
rect 422294 244876 422300 244888
rect 422352 244876 422358 244928
rect 73154 243516 73160 243568
rect 73212 243556 73218 243568
rect 273438 243556 273444 243568
rect 73212 243528 273444 243556
rect 73212 243516 73218 243528
rect 273438 243516 273444 243528
rect 273496 243516 273502 243568
rect 387886 243516 387892 243568
rect 387944 243556 387950 243568
rect 560294 243556 560300 243568
rect 387944 243528 560300 243556
rect 387944 243516 387950 243528
rect 560294 243516 560300 243528
rect 560352 243516 560358 243568
rect 80054 242156 80060 242208
rect 80112 242196 80118 242208
rect 274726 242196 274732 242208
rect 80112 242168 274732 242196
rect 80112 242156 80118 242168
rect 274726 242156 274732 242168
rect 274784 242156 274790 242208
rect 389358 242156 389364 242208
rect 389416 242196 389422 242208
rect 567194 242196 567200 242208
rect 389416 242168 567200 242196
rect 389416 242156 389422 242168
rect 567194 242156 567200 242168
rect 567252 242156 567258 242208
rect 3510 241408 3516 241460
rect 3568 241448 3574 241460
rect 220078 241448 220084 241460
rect 3568 241420 220084 241448
rect 3568 241408 3574 241420
rect 220078 241408 220084 241420
rect 220136 241408 220142 241460
rect 237466 240728 237472 240780
rect 237524 240768 237530 240780
rect 312170 240768 312176 240780
rect 237524 240740 312176 240768
rect 237524 240728 237530 240740
rect 312170 240728 312176 240740
rect 312228 240728 312234 240780
rect 393958 240728 393964 240780
rect 394016 240768 394022 240780
rect 578234 240768 578240 240780
rect 394016 240740 578240 240768
rect 394016 240728 394022 240740
rect 578234 240728 578240 240740
rect 578292 240728 578298 240780
rect 93946 239368 93952 239420
rect 94004 239408 94010 239420
rect 278866 239408 278872 239420
rect 94004 239380 278872 239408
rect 94004 239368 94010 239380
rect 278866 239368 278872 239380
rect 278924 239368 278930 239420
rect 111794 238008 111800 238060
rect 111852 238048 111858 238060
rect 283098 238048 283104 238060
rect 111852 238020 283104 238048
rect 111852 238008 111858 238020
rect 283098 238008 283104 238020
rect 283156 238008 283162 238060
rect 115934 236648 115940 236700
rect 115992 236688 115998 236700
rect 283006 236688 283012 236700
rect 115992 236660 283012 236688
rect 115992 236648 115998 236660
rect 283006 236648 283012 236660
rect 283064 236648 283070 236700
rect 30374 235220 30380 235272
rect 30432 235260 30438 235272
rect 263778 235260 263784 235272
rect 30432 235232 263784 235260
rect 30432 235220 30438 235232
rect 263778 235220 263784 235232
rect 263836 235220 263842 235272
rect 39298 233860 39304 233912
rect 39356 233900 39362 233912
rect 265158 233900 265164 233912
rect 39356 233872 265164 233900
rect 39356 233860 39362 233872
rect 265158 233860 265164 233872
rect 265216 233860 265222 233912
rect 395430 233180 395436 233232
rect 395488 233220 395494 233232
rect 580166 233220 580172 233232
rect 395488 233192 580172 233220
rect 395488 233180 395494 233192
rect 580166 233180 580172 233192
rect 580224 233180 580230 233232
rect 44266 232500 44272 232552
rect 44324 232540 44330 232552
rect 266446 232540 266452 232552
rect 44324 232512 266452 232540
rect 44324 232500 44330 232512
rect 266446 232500 266452 232512
rect 266504 232500 266510 232552
rect 49694 231072 49700 231124
rect 49752 231112 49758 231124
rect 267826 231112 267832 231124
rect 49752 231084 267832 231112
rect 49752 231072 49758 231084
rect 267826 231072 267832 231084
rect 267884 231072 267890 231124
rect 52546 229712 52552 229764
rect 52604 229752 52610 229764
rect 269298 229752 269304 229764
rect 52604 229724 269304 229752
rect 52604 229712 52610 229724
rect 269298 229712 269304 229724
rect 269356 229712 269362 229764
rect 56594 228352 56600 228404
rect 56652 228392 56658 228404
rect 269206 228392 269212 228404
rect 56652 228364 269212 228392
rect 56652 228352 56658 228364
rect 269206 228352 269212 228364
rect 269264 228352 269270 228404
rect 67634 226992 67640 227044
rect 67692 227032 67698 227044
rect 272150 227032 272156 227044
rect 67692 227004 272156 227032
rect 67692 226992 67698 227004
rect 272150 226992 272156 227004
rect 272208 226992 272214 227044
rect 74534 225564 74540 225616
rect 74592 225604 74598 225616
rect 273346 225604 273352 225616
rect 74592 225576 273352 225604
rect 74592 225564 74598 225576
rect 273346 225564 273352 225576
rect 273404 225564 273410 225616
rect 13814 224204 13820 224256
rect 13872 224244 13878 224256
rect 259638 224244 259644 224256
rect 13872 224216 259644 224244
rect 13872 224204 13878 224216
rect 259638 224204 259644 224216
rect 259696 224204 259702 224256
rect 158714 222844 158720 222896
rect 158772 222884 158778 222896
rect 293310 222884 293316 222896
rect 158772 222856 293316 222884
rect 158772 222844 158778 222856
rect 293310 222844 293316 222856
rect 293368 222844 293374 222896
rect 85666 221416 85672 221468
rect 85724 221456 85730 221468
rect 276290 221456 276296 221468
rect 85724 221428 276296 221456
rect 85724 221416 85730 221428
rect 276290 221416 276296 221428
rect 276348 221416 276354 221468
rect 92474 220056 92480 220108
rect 92532 220096 92538 220108
rect 277578 220096 277584 220108
rect 92532 220068 277584 220096
rect 92532 220056 92538 220068
rect 277578 220056 277584 220068
rect 277636 220056 277642 220108
rect 432598 219376 432604 219428
rect 432656 219416 432662 219428
rect 579890 219416 579896 219428
rect 432656 219388 579896 219416
rect 432656 219376 432662 219388
rect 579890 219376 579896 219388
rect 579948 219376 579954 219428
rect 102226 218696 102232 218748
rect 102284 218736 102290 218748
rect 280430 218736 280436 218748
rect 102284 218708 280436 218736
rect 102284 218696 102290 218708
rect 280430 218696 280436 218708
rect 280488 218696 280494 218748
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 18690 215268 18696 215280
rect 3384 215240 18696 215268
rect 3384 215228 3390 215240
rect 18690 215228 18696 215240
rect 18748 215228 18754 215280
rect 17954 214548 17960 214600
rect 18012 214588 18018 214600
rect 261018 214588 261024 214600
rect 18012 214560 261024 214588
rect 18012 214548 18018 214560
rect 261018 214548 261024 214560
rect 261076 214548 261082 214600
rect 421558 206932 421564 206984
rect 421616 206972 421622 206984
rect 580166 206972 580172 206984
rect 421616 206944 580172 206972
rect 421616 206932 421622 206944
rect 580166 206932 580172 206944
rect 580224 206932 580230 206984
rect 3050 202784 3056 202836
rect 3108 202824 3114 202836
rect 90358 202824 90364 202836
rect 3108 202796 90364 202824
rect 3108 202784 3114 202796
rect 90358 202784 90364 202796
rect 90416 202784 90422 202836
rect 428458 193128 428464 193180
rect 428516 193168 428522 193180
rect 580166 193168 580172 193180
rect 428516 193140 580172 193168
rect 428516 193128 428522 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 3510 188980 3516 189032
rect 3568 189020 3574 189032
rect 217318 189020 217324 189032
rect 3568 188992 217324 189020
rect 3568 188980 3574 188992
rect 217318 188980 217324 188992
rect 217376 188980 217382 189032
rect 216674 188300 216680 188352
rect 216732 188340 216738 188352
rect 306650 188340 306656 188352
rect 216732 188312 306656 188340
rect 216732 188300 216738 188312
rect 306650 188300 306656 188312
rect 306708 188300 306714 188352
rect 386506 182792 386512 182844
rect 386564 182832 386570 182844
rect 558914 182832 558920 182844
rect 386564 182804 558920 182832
rect 386564 182792 386570 182804
rect 558914 182792 558920 182804
rect 558972 182792 558978 182844
rect 404998 179324 405004 179376
rect 405056 179364 405062 179376
rect 579982 179364 579988 179376
rect 405056 179336 579988 179364
rect 405056 179324 405062 179336
rect 579982 179324 579988 179336
rect 580040 179324 580046 179376
rect 350626 178644 350632 178696
rect 350684 178684 350690 178696
rect 404354 178684 404360 178696
rect 350684 178656 404360 178684
rect 350684 178644 350690 178656
rect 404354 178644 404360 178656
rect 404412 178644 404418 178696
rect 390738 171776 390744 171828
rect 390796 171816 390802 171828
rect 574094 171816 574100 171828
rect 390796 171788 574100 171816
rect 390796 171776 390802 171788
rect 574094 171776 574100 171788
rect 574152 171776 574158 171828
rect 418798 166948 418804 167000
rect 418856 166988 418862 167000
rect 580166 166988 580172 167000
rect 418856 166960 580172 166988
rect 418856 166948 418862 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 251266 166268 251272 166320
rect 251324 166308 251330 166320
rect 314746 166308 314752 166320
rect 251324 166280 314752 166308
rect 251324 166268 251330 166280
rect 314746 166268 314752 166280
rect 314804 166268 314810 166320
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 229738 164200 229744 164212
rect 3292 164172 229744 164200
rect 3292 164160 3298 164172
rect 229738 164160 229744 164172
rect 229796 164160 229802 164212
rect 554038 153144 554044 153196
rect 554096 153184 554102 153196
rect 579798 153184 579804 153196
rect 554096 153156 579804 153184
rect 554096 153144 554102 153156
rect 579798 153144 579804 153156
rect 579856 153144 579862 153196
rect 346486 140020 346492 140072
rect 346544 140060 346550 140072
rect 386506 140060 386512 140072
rect 346544 140032 386512 140060
rect 346544 140020 346550 140032
rect 386506 140020 386512 140032
rect 386564 140020 386570 140072
rect 3510 137232 3516 137284
rect 3568 137272 3574 137284
rect 414106 137272 414112 137284
rect 3568 137244 414112 137272
rect 3568 137232 3574 137244
rect 414106 137232 414112 137244
rect 414164 137232 414170 137284
rect 417418 126896 417424 126948
rect 417476 126936 417482 126948
rect 580166 126936 580172 126948
rect 417476 126908 580172 126936
rect 417476 126896 417482 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 427078 113092 427084 113144
rect 427136 113132 427142 113144
rect 580166 113132 580172 113144
rect 427136 113104 580172 113132
rect 427136 113092 427142 113104
rect 580166 113092 580172 113104
rect 580224 113092 580230 113144
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 228358 111772 228364 111784
rect 3200 111744 228364 111772
rect 3200 111732 3206 111744
rect 228358 111732 228364 111744
rect 228416 111732 228422 111784
rect 250438 100648 250444 100700
rect 250496 100688 250502 100700
rect 580166 100688 580172 100700
rect 250496 100660 580172 100688
rect 250496 100648 250502 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 389266 90312 389272 90364
rect 389324 90352 389330 90364
rect 570598 90352 570604 90364
rect 389324 90324 570604 90352
rect 389324 90312 389330 90324
rect 570598 90312 570604 90324
rect 570656 90312 570662 90364
rect 414658 86912 414664 86964
rect 414716 86952 414722 86964
rect 580166 86952 580172 86964
rect 414716 86924 580172 86952
rect 414716 86912 414722 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 350534 86232 350540 86284
rect 350592 86272 350598 86284
rect 400214 86272 400220 86284
rect 350592 86244 400220 86272
rect 350592 86232 350598 86244
rect 400214 86232 400220 86244
rect 400272 86232 400278 86284
rect 3418 85484 3424 85536
rect 3476 85524 3482 85536
rect 400858 85524 400864 85536
rect 3476 85496 400864 85524
rect 3476 85484 3482 85496
rect 400858 85484 400864 85496
rect 400916 85484 400922 85536
rect 424318 73108 424324 73160
rect 424376 73148 424382 73160
rect 579982 73148 579988 73160
rect 424376 73120 579988 73148
rect 424376 73108 424382 73120
rect 579982 73108 579988 73120
rect 580040 73108 580046 73160
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 225598 71720 225604 71732
rect 3476 71692 225604 71720
rect 3476 71680 3482 71692
rect 225598 71680 225604 71692
rect 225656 71680 225662 71732
rect 246298 60664 246304 60716
rect 246356 60704 246362 60716
rect 580166 60704 580172 60716
rect 246356 60676 580172 60704
rect 246356 60664 246362 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 127066 51688 127072 51740
rect 127124 51728 127130 51740
rect 285858 51728 285864 51740
rect 127124 51700 285864 51728
rect 127124 51688 127130 51700
rect 285858 51688 285864 51700
rect 285916 51688 285922 51740
rect 285950 51688 285956 51740
rect 286008 51728 286014 51740
rect 323118 51728 323124 51740
rect 286008 51700 323124 51728
rect 286008 51688 286014 51700
rect 323118 51688 323124 51700
rect 323176 51688 323182 51740
rect 113174 48968 113180 49020
rect 113232 49008 113238 49020
rect 282914 49008 282920 49020
rect 113232 48980 282920 49008
rect 113232 48968 113238 48980
rect 282914 48968 282920 48980
rect 282972 48968 282978 49020
rect 345198 47676 345204 47728
rect 345256 47716 345262 47728
rect 382550 47716 382556 47728
rect 345256 47688 382556 47716
rect 345256 47676 345262 47688
rect 382550 47676 382556 47688
rect 382608 47676 382614 47728
rect 95234 47540 95240 47592
rect 95292 47580 95298 47592
rect 279142 47580 279148 47592
rect 95292 47552 279148 47580
rect 95292 47540 95298 47552
rect 279142 47540 279148 47552
rect 279200 47540 279206 47592
rect 382366 47540 382372 47592
rect 382424 47580 382430 47592
rect 540974 47580 540980 47592
rect 382424 47552 540980 47580
rect 382424 47540 382430 47552
rect 540974 47540 540980 47552
rect 541032 47540 541038 47592
rect 238018 46180 238024 46232
rect 238076 46220 238082 46232
rect 580350 46220 580356 46232
rect 238076 46192 580356 46220
rect 238076 46180 238082 46192
rect 580350 46180 580356 46192
rect 580408 46180 580414 46232
rect 122834 43392 122840 43444
rect 122892 43432 122898 43444
rect 285766 43432 285772 43444
rect 122892 43404 285772 43432
rect 122892 43392 122898 43404
rect 285766 43392 285772 43404
rect 285824 43392 285830 43444
rect 77386 42032 77392 42084
rect 77444 42072 77450 42084
rect 275002 42072 275008 42084
rect 77444 42044 275008 42072
rect 77444 42032 77450 42044
rect 275002 42032 275008 42044
rect 275060 42032 275066 42084
rect 9674 40672 9680 40724
rect 9732 40712 9738 40724
rect 257430 40712 257436 40724
rect 9732 40684 257436 40712
rect 9732 40672 9738 40684
rect 257430 40672 257436 40684
rect 257488 40672 257494 40724
rect 69106 39312 69112 39364
rect 69164 39352 69170 39364
rect 271138 39352 271144 39364
rect 69164 39324 271144 39352
rect 69164 39312 69170 39324
rect 271138 39312 271144 39324
rect 271196 39312 271202 39364
rect 140774 37884 140780 37936
rect 140832 37924 140838 37936
rect 289078 37924 289084 37936
rect 140832 37896 289084 37924
rect 140832 37884 140838 37896
rect 289078 37884 289084 37896
rect 289136 37884 289142 37936
rect 55214 36524 55220 36576
rect 55272 36564 55278 36576
rect 269482 36564 269488 36576
rect 55272 36536 269488 36564
rect 55272 36524 55278 36536
rect 269482 36524 269488 36536
rect 269540 36524 269546 36576
rect 160186 35164 160192 35216
rect 160244 35204 160250 35216
rect 293218 35204 293224 35216
rect 160244 35176 293224 35204
rect 160244 35164 160250 35176
rect 293218 35164 293224 35176
rect 293276 35164 293282 35216
rect 244274 33736 244280 33788
rect 244332 33776 244338 33788
rect 313642 33776 313648 33788
rect 244332 33748 313648 33776
rect 244332 33736 244338 33748
rect 313642 33736 313648 33748
rect 313700 33736 313706 33788
rect 3418 33056 3424 33108
rect 3476 33096 3482 33108
rect 224218 33096 224224 33108
rect 3476 33068 224224 33096
rect 3476 33056 3482 33068
rect 224218 33056 224224 33068
rect 224276 33056 224282 33108
rect 237374 33056 237380 33108
rect 237432 33096 237438 33108
rect 580166 33096 580172 33108
rect 237432 33068 580172 33096
rect 237432 33056 237438 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 226426 31016 226432 31068
rect 226484 31056 226490 31068
rect 309502 31056 309508 31068
rect 226484 31028 309508 31056
rect 226484 31016 226490 31028
rect 309502 31016 309508 31028
rect 309560 31016 309566 31068
rect 212534 29588 212540 29640
rect 212592 29628 212598 29640
rect 302878 29628 302884 29640
rect 212592 29600 302884 29628
rect 212592 29588 212598 29600
rect 302878 29588 302884 29600
rect 302936 29588 302942 29640
rect 352006 29588 352012 29640
rect 352064 29628 352070 29640
rect 407206 29628 407212 29640
rect 352064 29600 407212 29628
rect 352064 29588 352070 29600
rect 407206 29588 407212 29600
rect 407264 29588 407270 29640
rect 209866 28228 209872 28280
rect 209924 28268 209930 28280
rect 305270 28268 305276 28280
rect 209924 28240 305276 28268
rect 209924 28228 209930 28240
rect 305270 28228 305276 28240
rect 305328 28228 305334 28280
rect 349338 28228 349344 28280
rect 349396 28268 349402 28280
rect 397454 28268 397460 28280
rect 349396 28240 397460 28268
rect 349396 28228 349402 28240
rect 397454 28228 397460 28240
rect 397512 28228 397518 28280
rect 194594 26868 194600 26920
rect 194652 26908 194658 26920
rect 302234 26908 302240 26920
rect 194652 26880 302240 26908
rect 194652 26868 194658 26880
rect 302234 26868 302240 26880
rect 302292 26868 302298 26920
rect 347774 26868 347780 26920
rect 347832 26908 347838 26920
rect 393314 26908 393320 26920
rect 347832 26880 393320 26908
rect 347832 26868 347838 26880
rect 393314 26868 393320 26880
rect 393372 26868 393378 26920
rect 186314 25508 186320 25560
rect 186372 25548 186378 25560
rect 299842 25548 299848 25560
rect 186372 25520 299848 25548
rect 186372 25508 186378 25520
rect 299842 25508 299848 25520
rect 299900 25508 299906 25560
rect 343634 25508 343640 25560
rect 343692 25548 343698 25560
rect 375374 25548 375380 25560
rect 343692 25520 375380 25548
rect 343692 25508 343698 25520
rect 375374 25508 375380 25520
rect 375432 25508 375438 25560
rect 176746 24080 176752 24132
rect 176804 24120 176810 24132
rect 296162 24120 296168 24132
rect 176804 24092 296168 24120
rect 176804 24080 176810 24092
rect 296162 24080 296168 24092
rect 296220 24080 296226 24132
rect 341058 24080 341064 24132
rect 341116 24120 341122 24132
rect 361574 24120 361580 24132
rect 341116 24092 361580 24120
rect 341116 24080 341122 24092
rect 361574 24080 361580 24092
rect 361632 24080 361638 24132
rect 382274 24080 382280 24132
rect 382332 24120 382338 24132
rect 539686 24120 539692 24132
rect 382332 24092 539692 24120
rect 382332 24080 382338 24092
rect 539686 24080 539692 24092
rect 539744 24080 539750 24132
rect 154574 22720 154580 22772
rect 154632 22760 154638 22772
rect 291838 22760 291844 22772
rect 154632 22732 291844 22760
rect 154632 22720 154638 22732
rect 291838 22720 291844 22732
rect 291896 22720 291902 22772
rect 292574 22720 292580 22772
rect 292632 22760 292638 22772
rect 324498 22760 324504 22772
rect 292632 22732 324504 22760
rect 292632 22720 292638 22732
rect 324498 22720 324504 22732
rect 324556 22720 324562 22772
rect 342438 22720 342444 22772
rect 342496 22760 342502 22772
rect 368658 22760 368664 22772
rect 342496 22732 368664 22760
rect 342496 22720 342502 22732
rect 368658 22720 368664 22732
rect 368716 22720 368722 22772
rect 380894 22720 380900 22772
rect 380952 22760 380958 22772
rect 531406 22760 531412 22772
rect 380952 22732 531412 22760
rect 380952 22720 380958 22732
rect 531406 22720 531412 22732
rect 531464 22720 531470 22772
rect 204254 21360 204260 21412
rect 204312 21400 204318 21412
rect 303706 21400 303712 21412
rect 204312 21372 303712 21400
rect 204312 21360 204318 21372
rect 303706 21360 303712 21372
rect 303764 21360 303770 21412
rect 310514 21360 310520 21412
rect 310572 21400 310578 21412
rect 328730 21400 328736 21412
rect 310572 21372 328736 21400
rect 310572 21360 310578 21372
rect 328730 21360 328736 21372
rect 328788 21360 328794 21412
rect 337102 21360 337108 21412
rect 337160 21400 337166 21412
rect 346486 21400 346492 21412
rect 337160 21372 346492 21400
rect 337160 21360 337166 21372
rect 346486 21360 346492 21372
rect 346544 21360 346550 21412
rect 376754 21360 376760 21412
rect 376812 21400 376818 21412
rect 514754 21400 514760 21412
rect 376812 21372 514760 21400
rect 376812 21360 376818 21372
rect 514754 21360 514760 21372
rect 514812 21360 514818 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 413370 20652 413376 20664
rect 3476 20624 413376 20652
rect 3476 20612 3482 20624
rect 413370 20612 413376 20624
rect 413428 20612 413434 20664
rect 269114 18640 269120 18692
rect 269172 18680 269178 18692
rect 319070 18680 319076 18692
rect 269172 18652 319076 18680
rect 269172 18640 269178 18652
rect 319070 18640 319076 18652
rect 319128 18640 319134 18692
rect 172514 18572 172520 18624
rect 172572 18612 172578 18624
rect 296070 18612 296076 18624
rect 172572 18584 296076 18612
rect 172572 18572 172578 18584
rect 296070 18572 296076 18584
rect 296128 18572 296134 18624
rect 299474 18572 299480 18624
rect 299532 18612 299538 18624
rect 323670 18612 323676 18624
rect 299532 18584 323676 18612
rect 299532 18572 299538 18584
rect 323670 18572 323676 18584
rect 323728 18572 323734 18624
rect 368566 18572 368572 18624
rect 368624 18612 368630 18624
rect 481726 18612 481732 18624
rect 368624 18584 481732 18612
rect 368624 18572 368630 18584
rect 481726 18572 481732 18584
rect 481784 18572 481790 18624
rect 259638 17280 259644 17332
rect 259696 17320 259702 17332
rect 317598 17320 317604 17332
rect 259696 17292 317604 17320
rect 259696 17280 259702 17292
rect 317598 17280 317604 17292
rect 317656 17280 317662 17332
rect 349154 17280 349160 17332
rect 349212 17320 349218 17332
rect 398926 17320 398932 17332
rect 349212 17292 398932 17320
rect 349212 17280 349218 17292
rect 398926 17280 398932 17292
rect 398984 17280 398990 17332
rect 118786 17212 118792 17264
rect 118844 17252 118850 17264
rect 284478 17252 284484 17264
rect 118844 17224 284484 17252
rect 118844 17212 118850 17224
rect 284478 17212 284484 17224
rect 284536 17212 284542 17264
rect 295334 17212 295340 17264
rect 295392 17252 295398 17264
rect 324958 17252 324964 17264
rect 295392 17224 324964 17252
rect 295392 17212 295398 17224
rect 324958 17212 324964 17224
rect 325016 17212 325022 17264
rect 387794 17212 387800 17264
rect 387852 17252 387858 17264
rect 564526 17252 564532 17264
rect 387852 17224 564532 17252
rect 387852 17212 387858 17224
rect 564526 17212 564532 17224
rect 564584 17212 564590 17264
rect 109034 16056 109040 16108
rect 109092 16096 109098 16108
rect 281626 16096 281632 16108
rect 109092 16068 281632 16096
rect 109092 16056 109098 16068
rect 281626 16056 281632 16068
rect 281684 16056 281690 16108
rect 105722 15988 105728 16040
rect 105780 16028 105786 16040
rect 281718 16028 281724 16040
rect 105780 16000 281724 16028
rect 105780 15988 105786 16000
rect 281718 15988 281724 16000
rect 281776 15988 281782 16040
rect 91554 15920 91560 15972
rect 91612 15960 91618 15972
rect 277394 15960 277400 15972
rect 91612 15932 277400 15960
rect 91612 15920 91618 15932
rect 277394 15920 277400 15932
rect 277452 15920 277458 15972
rect 281994 15920 282000 15972
rect 282052 15960 282058 15972
rect 304258 15960 304264 15972
rect 282052 15932 304264 15960
rect 282052 15920 282058 15932
rect 304258 15920 304264 15932
rect 304316 15920 304322 15972
rect 345106 15920 345112 15972
rect 345164 15960 345170 15972
rect 379514 15960 379520 15972
rect 345164 15932 379520 15960
rect 345164 15920 345170 15932
rect 379514 15920 379520 15932
rect 379572 15920 379578 15972
rect 87506 15852 87512 15904
rect 87564 15892 87570 15904
rect 277486 15892 277492 15904
rect 87564 15864 277492 15892
rect 87564 15852 87570 15864
rect 277486 15852 277492 15864
rect 277544 15852 277550 15904
rect 279050 15852 279056 15904
rect 279108 15892 279114 15904
rect 316678 15892 316684 15904
rect 279108 15864 316684 15892
rect 279108 15852 279114 15864
rect 316678 15852 316684 15864
rect 316736 15852 316742 15904
rect 372614 15852 372620 15904
rect 372672 15892 372678 15904
rect 497090 15892 497096 15904
rect 372672 15864 497096 15892
rect 372672 15852 372678 15864
rect 497090 15852 497096 15864
rect 497148 15852 497154 15904
rect 273346 14560 273352 14612
rect 273404 14600 273410 14612
rect 320358 14600 320364 14612
rect 273404 14572 320364 14600
rect 273404 14560 273410 14572
rect 320358 14560 320364 14572
rect 320416 14560 320422 14612
rect 122282 14492 122288 14544
rect 122340 14532 122346 14544
rect 284386 14532 284392 14544
rect 122340 14504 284392 14532
rect 122340 14492 122346 14504
rect 284386 14492 284392 14504
rect 284444 14492 284450 14544
rect 108114 14424 108120 14476
rect 108172 14464 108178 14476
rect 281902 14464 281908 14476
rect 108172 14436 281908 14464
rect 108172 14424 108178 14436
rect 281902 14424 281908 14436
rect 281960 14424 281966 14476
rect 284570 14424 284576 14476
rect 284628 14464 284634 14476
rect 305638 14464 305644 14476
rect 284628 14436 305644 14464
rect 284628 14424 284634 14436
rect 305638 14424 305644 14436
rect 305696 14424 305702 14476
rect 306374 14424 306380 14476
rect 306432 14464 306438 14476
rect 328638 14464 328644 14476
rect 306432 14436 328644 14464
rect 306432 14424 306438 14436
rect 328638 14424 328644 14436
rect 328696 14424 328702 14476
rect 339586 14424 339592 14476
rect 339644 14464 339650 14476
rect 357526 14464 357532 14476
rect 339644 14436 357532 14464
rect 339644 14424 339650 14436
rect 357526 14424 357532 14436
rect 357584 14424 357590 14476
rect 378134 14424 378140 14476
rect 378192 14464 378198 14476
rect 523770 14464 523776 14476
rect 378192 14436 523776 14464
rect 378192 14424 378198 14436
rect 523770 14424 523776 14436
rect 523828 14424 523834 14476
rect 278314 13200 278320 13252
rect 278372 13240 278378 13252
rect 300118 13240 300124 13252
rect 278372 13212 300124 13240
rect 278372 13200 278378 13212
rect 300118 13200 300124 13212
rect 300176 13200 300182 13252
rect 283098 13132 283104 13184
rect 283156 13172 283162 13184
rect 307018 13172 307024 13184
rect 283156 13144 307024 13172
rect 283156 13132 283162 13144
rect 307018 13132 307024 13144
rect 307076 13132 307082 13184
rect 346394 13132 346400 13184
rect 346452 13172 346458 13184
rect 387794 13172 387800 13184
rect 346452 13144 387800 13172
rect 346452 13132 346458 13144
rect 387794 13132 387800 13144
rect 387852 13132 387858 13184
rect 137186 13064 137192 13116
rect 137244 13104 137250 13116
rect 287698 13104 287704 13116
rect 137244 13076 287704 13104
rect 137244 13064 137250 13076
rect 287698 13064 287704 13076
rect 287756 13064 287762 13116
rect 303154 13064 303160 13116
rect 303212 13104 303218 13116
rect 327258 13104 327264 13116
rect 303212 13076 327264 13104
rect 303212 13064 303218 13076
rect 327258 13064 327264 13076
rect 327316 13064 327322 13116
rect 386414 13064 386420 13116
rect 386472 13104 386478 13116
rect 556890 13104 556896 13116
rect 386472 13076 556896 13104
rect 386472 13064 386478 13076
rect 556890 13064 556896 13076
rect 556948 13064 556954 13116
rect 143534 11772 143540 11824
rect 143592 11812 143598 11824
rect 144730 11812 144736 11824
rect 143592 11784 144736 11812
rect 143592 11772 143598 11784
rect 144730 11772 144736 11784
rect 144788 11772 144794 11824
rect 160094 11772 160100 11824
rect 160152 11812 160158 11824
rect 161290 11812 161296 11824
rect 160152 11784 161296 11812
rect 160152 11772 160158 11784
rect 161290 11772 161296 11784
rect 161348 11772 161354 11824
rect 184934 11772 184940 11824
rect 184992 11812 184998 11824
rect 186130 11812 186136 11824
rect 184992 11784 186136 11812
rect 184992 11772 184998 11784
rect 186130 11772 186136 11784
rect 186188 11772 186194 11824
rect 234614 11772 234620 11824
rect 234672 11812 234678 11824
rect 235810 11812 235816 11824
rect 234672 11784 235816 11812
rect 234672 11772 234678 11784
rect 235810 11772 235816 11784
rect 235868 11772 235874 11824
rect 242894 11772 242900 11824
rect 242952 11812 242958 11824
rect 244090 11812 244096 11824
rect 242952 11784 244096 11812
rect 242952 11772 242958 11784
rect 244090 11772 244096 11784
rect 244148 11772 244154 11824
rect 274818 11772 274824 11824
rect 274876 11812 274882 11824
rect 320266 11812 320272 11824
rect 274876 11784 320272 11812
rect 274876 11772 274882 11784
rect 320266 11772 320272 11784
rect 320324 11772 320330 11824
rect 351914 11772 351920 11824
rect 351972 11812 351978 11824
rect 411898 11812 411904 11824
rect 351972 11784 411904 11812
rect 351972 11772 351978 11784
rect 411898 11772 411904 11784
rect 411956 11772 411962 11824
rect 51074 11704 51080 11756
rect 51132 11744 51138 11756
rect 257338 11744 257344 11756
rect 51132 11716 257344 11744
rect 51132 11704 51138 11716
rect 257338 11704 257344 11716
rect 257396 11704 257402 11756
rect 265158 11704 265164 11756
rect 265216 11744 265222 11756
rect 318978 11744 318984 11756
rect 265216 11716 318984 11744
rect 265216 11704 265222 11716
rect 318978 11704 318984 11716
rect 319036 11704 319042 11756
rect 340966 11704 340972 11756
rect 341024 11744 341030 11756
rect 363506 11744 363512 11756
rect 341024 11716 363512 11744
rect 341024 11704 341030 11716
rect 363506 11704 363512 11716
rect 363564 11704 363570 11756
rect 407758 11704 407764 11756
rect 407816 11744 407822 11756
rect 537202 11744 537208 11756
rect 407816 11716 537208 11744
rect 407816 11704 407822 11716
rect 537202 11704 537208 11716
rect 537260 11704 537266 11756
rect 309870 10480 309876 10532
rect 309928 10520 309934 10532
rect 328546 10520 328552 10532
rect 309928 10492 328552 10520
rect 309928 10480 309934 10492
rect 328546 10480 328552 10492
rect 328604 10480 328610 10532
rect 270770 10412 270776 10464
rect 270828 10452 270834 10464
rect 309778 10452 309784 10464
rect 270828 10424 309784 10452
rect 270828 10412 270834 10424
rect 309778 10412 309784 10424
rect 309836 10412 309842 10464
rect 280706 10344 280712 10396
rect 280764 10384 280770 10396
rect 321646 10384 321652 10396
rect 280764 10356 321652 10384
rect 280764 10344 280770 10356
rect 321646 10344 321652 10356
rect 321704 10344 321710 10396
rect 72602 10276 72608 10328
rect 72660 10316 72666 10328
rect 273622 10316 273628 10328
rect 72660 10288 273628 10316
rect 72660 10276 72666 10288
rect 273622 10276 273628 10288
rect 273680 10276 273686 10328
rect 276014 10276 276020 10328
rect 276072 10316 276078 10328
rect 320450 10316 320456 10328
rect 276072 10288 320456 10316
rect 276072 10276 276078 10288
rect 320450 10276 320456 10288
rect 320508 10276 320514 10328
rect 342346 10276 342352 10328
rect 342404 10316 342410 10328
rect 370130 10316 370136 10328
rect 342404 10288 370136 10316
rect 342404 10276 342410 10288
rect 370130 10276 370136 10288
rect 370188 10276 370194 10328
rect 399478 10276 399484 10328
rect 399536 10316 399542 10328
rect 515490 10316 515496 10328
rect 399536 10288 515496 10316
rect 399536 10276 399542 10288
rect 515490 10276 515496 10288
rect 515548 10276 515554 10328
rect 209682 9596 209688 9648
rect 209740 9636 209746 9648
rect 210970 9636 210976 9648
rect 209740 9608 210976 9636
rect 209740 9596 209746 9608
rect 210970 9596 210976 9608
rect 211028 9596 211034 9648
rect 359458 9596 359464 9648
rect 359516 9636 359522 9648
rect 361114 9636 361120 9648
rect 359516 9608 361120 9636
rect 359516 9596 359522 9608
rect 361114 9596 361120 9608
rect 361172 9596 361178 9648
rect 261754 9052 261760 9104
rect 261812 9092 261818 9104
rect 311158 9092 311164 9104
rect 261812 9064 311164 9092
rect 261812 9052 261818 9064
rect 311158 9052 311164 9064
rect 311216 9052 311222 9104
rect 266538 8984 266544 9036
rect 266596 9024 266602 9036
rect 318886 9024 318892 9036
rect 266596 8996 318892 9024
rect 266596 8984 266602 8996
rect 318886 8984 318892 8996
rect 318944 8984 318950 9036
rect 132954 8916 132960 8968
rect 133012 8956 133018 8968
rect 243538 8956 243544 8968
rect 133012 8928 243544 8956
rect 133012 8916 133018 8928
rect 243538 8916 243544 8928
rect 243596 8916 243602 8968
rect 264146 8916 264152 8968
rect 264204 8956 264210 8968
rect 317506 8956 317512 8968
rect 264204 8928 317512 8956
rect 264204 8916 264210 8928
rect 317506 8916 317512 8928
rect 317564 8916 317570 8968
rect 320910 8916 320916 8968
rect 320968 8956 320974 8968
rect 331490 8956 331496 8968
rect 320968 8928 331496 8956
rect 320968 8916 320974 8928
rect 331490 8916 331496 8928
rect 331548 8916 331554 8968
rect 340874 8916 340880 8968
rect 340932 8956 340938 8968
rect 359918 8956 359924 8968
rect 340932 8928 359924 8956
rect 340932 8916 340938 8928
rect 359918 8916 359924 8928
rect 359976 8916 359982 8968
rect 370498 8916 370504 8968
rect 370556 8956 370562 8968
rect 393038 8956 393044 8968
rect 370556 8928 393044 8956
rect 370556 8916 370562 8928
rect 393038 8916 393044 8928
rect 393096 8916 393102 8968
rect 410518 8916 410524 8968
rect 410576 8956 410582 8968
rect 501782 8956 501788 8968
rect 410576 8928 501788 8956
rect 410576 8916 410582 8928
rect 501782 8916 501788 8928
rect 501840 8916 501846 8968
rect 360838 8372 360844 8424
rect 360896 8412 360902 8424
rect 365806 8412 365812 8424
rect 360896 8384 365812 8412
rect 360896 8372 360902 8384
rect 365806 8372 365812 8384
rect 365864 8372 365870 8424
rect 292574 7760 292580 7812
rect 292632 7800 292638 7812
rect 324406 7800 324412 7812
rect 292632 7772 324412 7800
rect 292632 7760 292638 7772
rect 324406 7760 324412 7772
rect 324464 7760 324470 7812
rect 260650 7692 260656 7744
rect 260708 7732 260714 7744
rect 301498 7732 301504 7744
rect 260708 7704 301504 7732
rect 260708 7692 260714 7704
rect 301498 7692 301504 7704
rect 301556 7692 301562 7744
rect 218146 7624 218152 7676
rect 218204 7664 218210 7676
rect 247678 7664 247684 7676
rect 218204 7636 247684 7664
rect 218204 7624 218210 7636
rect 247678 7624 247684 7636
rect 247736 7624 247742 7676
rect 277118 7624 277124 7676
rect 277176 7664 277182 7676
rect 321738 7664 321744 7676
rect 277176 7636 321744 7664
rect 277176 7624 277182 7636
rect 321738 7624 321744 7636
rect 321796 7624 321802 7676
rect 338390 7624 338396 7676
rect 338448 7664 338454 7676
rect 349154 7664 349160 7676
rect 338448 7636 349160 7664
rect 338448 7624 338454 7636
rect 349154 7624 349160 7636
rect 349212 7624 349218 7676
rect 33594 7556 33600 7608
rect 33652 7596 33658 7608
rect 233878 7596 233884 7608
rect 33652 7568 233884 7596
rect 33652 7556 33658 7568
rect 233878 7556 233884 7568
rect 233936 7556 233942 7608
rect 268838 7556 268844 7608
rect 268896 7596 268902 7608
rect 319162 7596 319168 7608
rect 268896 7568 319168 7596
rect 268896 7556 268902 7568
rect 319162 7556 319168 7568
rect 319220 7556 319226 7608
rect 324406 7556 324412 7608
rect 324464 7596 324470 7608
rect 332962 7596 332968 7608
rect 324464 7568 332968 7596
rect 324464 7556 324470 7568
rect 332962 7556 332968 7568
rect 333020 7556 333026 7608
rect 345014 7556 345020 7608
rect 345072 7596 345078 7608
rect 381170 7596 381176 7608
rect 345072 7568 381176 7596
rect 345072 7556 345078 7568
rect 381170 7556 381176 7568
rect 381228 7556 381234 7608
rect 395338 7556 395344 7608
rect 395396 7596 395402 7608
rect 487614 7596 487620 7608
rect 395396 7568 487620 7596
rect 395396 7556 395402 7568
rect 487614 7556 487620 7568
rect 487672 7556 487678 7608
rect 235994 6808 236000 6860
rect 236052 6848 236058 6860
rect 580166 6848 580172 6860
rect 236052 6820 580172 6848
rect 236052 6808 236058 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 288986 6264 288992 6316
rect 289044 6304 289050 6316
rect 297358 6304 297364 6316
rect 289044 6276 297364 6304
rect 289044 6264 289050 6276
rect 297358 6264 297364 6276
rect 297416 6264 297422 6316
rect 262950 6196 262956 6248
rect 263008 6236 263014 6248
rect 317690 6236 317696 6248
rect 263008 6208 317696 6236
rect 263008 6196 263014 6208
rect 317690 6196 317696 6208
rect 317748 6196 317754 6248
rect 169570 6128 169576 6180
rect 169628 6168 169634 6180
rect 242158 6168 242164 6180
rect 169628 6140 242164 6168
rect 169628 6128 169634 6140
rect 242158 6128 242164 6140
rect 242216 6128 242222 6180
rect 258258 6128 258264 6180
rect 258316 6168 258322 6180
rect 315298 6168 315304 6180
rect 258316 6140 315304 6168
rect 258316 6128 258322 6140
rect 315298 6128 315304 6140
rect 315356 6128 315362 6180
rect 318518 6128 318524 6180
rect 318576 6168 318582 6180
rect 327718 6168 327724 6180
rect 318576 6140 327724 6168
rect 318576 6128 318582 6140
rect 327718 6128 327724 6140
rect 327776 6128 327782 6180
rect 339494 6128 339500 6180
rect 339552 6168 339558 6180
rect 358722 6168 358728 6180
rect 339552 6140 358728 6168
rect 339552 6128 339558 6140
rect 358722 6128 358728 6140
rect 358780 6128 358786 6180
rect 267734 4972 267740 5024
rect 267792 5012 267798 5024
rect 295978 5012 295984 5024
rect 267792 4984 295984 5012
rect 267792 4972 267798 4984
rect 295978 4972 295984 4984
rect 296036 4972 296042 5024
rect 313826 4972 313832 5024
rect 313884 5012 313890 5024
rect 320818 5012 320824 5024
rect 313884 4984 320824 5012
rect 313884 4972 313890 4984
rect 320818 4972 320824 4984
rect 320876 4972 320882 5024
rect 290182 4904 290188 4956
rect 290240 4944 290246 4956
rect 323578 4944 323584 4956
rect 290240 4916 323584 4944
rect 290240 4904 290246 4916
rect 323578 4904 323584 4916
rect 323636 4904 323642 4956
rect 336918 4904 336924 4956
rect 336976 4944 336982 4956
rect 345750 4944 345756 4956
rect 336976 4916 345756 4944
rect 336976 4904 336982 4916
rect 345750 4904 345756 4916
rect 345808 4904 345814 4956
rect 272426 4836 272432 4888
rect 272484 4876 272490 4888
rect 318058 4876 318064 4888
rect 272484 4848 318064 4876
rect 272484 4836 272490 4848
rect 318058 4836 318064 4848
rect 318116 4836 318122 4888
rect 338298 4836 338304 4888
rect 338356 4876 338362 4888
rect 352834 4876 352840 4888
rect 338356 4848 352840 4876
rect 338356 4836 338362 4848
rect 352834 4836 352840 4848
rect 352892 4836 352898 4888
rect 353294 4836 353300 4888
rect 353352 4876 353358 4888
rect 415486 4876 415492 4888
rect 353352 4848 415492 4876
rect 353352 4836 353358 4848
rect 415486 4836 415492 4848
rect 415544 4836 415550 4888
rect 168374 4768 168380 4820
rect 168432 4808 168438 4820
rect 255958 4808 255964 4820
rect 168432 4780 255964 4808
rect 168432 4768 168438 4780
rect 255958 4768 255964 4780
rect 256016 4768 256022 4820
rect 257062 4768 257068 4820
rect 257120 4808 257126 4820
rect 313918 4808 313924 4820
rect 257120 4780 313924 4808
rect 257120 4768 257126 4780
rect 313918 4768 313924 4780
rect 313976 4768 313982 4820
rect 342254 4768 342260 4820
rect 342312 4808 342318 4820
rect 342312 4780 354674 4808
rect 342312 4768 342318 4780
rect 354646 4740 354674 4780
rect 363598 4768 363604 4820
rect 363656 4808 363662 4820
rect 364610 4808 364616 4820
rect 363656 4780 364616 4808
rect 363656 4768 363662 4780
rect 364610 4768 364616 4780
rect 364668 4768 364674 4820
rect 371878 4768 371884 4820
rect 371936 4808 371942 4820
rect 377674 4808 377680 4820
rect 371936 4780 377680 4808
rect 371936 4768 371942 4780
rect 377674 4768 377680 4780
rect 377732 4768 377738 4820
rect 396718 4768 396724 4820
rect 396776 4808 396782 4820
rect 484026 4808 484032 4820
rect 396776 4780 484032 4808
rect 396776 4768 396782 4780
rect 484026 4768 484032 4780
rect 484084 4768 484090 4820
rect 367002 4740 367008 4752
rect 354646 4712 367008 4740
rect 367002 4700 367008 4712
rect 367060 4700 367066 4752
rect 378778 4496 378784 4548
rect 378836 4536 378842 4548
rect 384758 4536 384764 4548
rect 378836 4508 384764 4536
rect 378836 4496 378842 4508
rect 384758 4496 384764 4508
rect 384816 4496 384822 4548
rect 135254 4156 135260 4208
rect 135312 4196 135318 4208
rect 136450 4196 136456 4208
rect 135312 4168 136456 4196
rect 135312 4156 135318 4168
rect 136450 4156 136456 4168
rect 136508 4156 136514 4208
rect 218054 4156 218060 4208
rect 218112 4196 218118 4208
rect 219250 4196 219256 4208
rect 218112 4168 219256 4196
rect 218112 4156 218118 4168
rect 219250 4156 219256 4168
rect 219308 4156 219314 4208
rect 258442 4196 258448 4208
rect 258276 4168 258448 4196
rect 43070 4088 43076 4140
rect 43128 4128 43134 4140
rect 258276 4128 258304 4168
rect 258442 4156 258448 4168
rect 258500 4156 258506 4208
rect 317322 4156 317328 4208
rect 317380 4196 317386 4208
rect 322198 4196 322204 4208
rect 317380 4168 322204 4196
rect 317380 4156 317386 4168
rect 322198 4156 322204 4168
rect 322256 4156 322262 4208
rect 337010 4156 337016 4208
rect 337068 4196 337074 4208
rect 342162 4196 342168 4208
rect 337068 4168 342168 4196
rect 337068 4156 337074 4168
rect 342162 4156 342168 4168
rect 342220 4156 342226 4208
rect 43128 4100 258304 4128
rect 43128 4088 43134 4100
rect 319714 4088 319720 4140
rect 319772 4128 319778 4140
rect 331398 4128 331404 4140
rect 319772 4100 331404 4128
rect 319772 4088 319778 4100
rect 331398 4088 331404 4100
rect 331456 4088 331462 4140
rect 358814 4088 358820 4140
rect 358872 4128 358878 4140
rect 440234 4128 440240 4140
rect 358872 4100 440240 4128
rect 358872 4088 358878 4100
rect 440234 4088 440240 4100
rect 440292 4088 440298 4140
rect 2866 4020 2872 4072
rect 2924 4060 2930 4072
rect 8938 4060 8944 4072
rect 2924 4032 8944 4060
rect 2924 4020 2930 4032
rect 8938 4020 8944 4032
rect 8996 4020 9002 4072
rect 39574 4020 39580 4072
rect 39632 4060 39638 4072
rect 265066 4060 265072 4072
rect 39632 4032 265072 4060
rect 39632 4020 39638 4032
rect 265066 4020 265072 4032
rect 265124 4020 265130 4072
rect 316218 4020 316224 4072
rect 316276 4060 316282 4072
rect 330110 4060 330116 4072
rect 316276 4032 330116 4060
rect 316276 4020 316282 4032
rect 330110 4020 330116 4032
rect 330168 4020 330174 4072
rect 360194 4020 360200 4072
rect 360252 4060 360258 4072
rect 447410 4060 447416 4072
rect 360252 4032 447416 4060
rect 360252 4020 360258 4032
rect 447410 4020 447416 4032
rect 447468 4020 447474 4072
rect 35986 3952 35992 4004
rect 36044 3992 36050 4004
rect 264974 3992 264980 4004
rect 36044 3964 264980 3992
rect 36044 3952 36050 3964
rect 264974 3952 264980 3964
rect 265032 3952 265038 4004
rect 312630 3952 312636 4004
rect 312688 3992 312694 4004
rect 329926 3992 329932 4004
rect 312688 3964 329932 3992
rect 312688 3952 312694 3964
rect 329926 3952 329932 3964
rect 329984 3952 329990 4004
rect 362954 3952 362960 4004
rect 363012 3992 363018 4004
rect 454494 3992 454500 4004
rect 363012 3964 454500 3992
rect 363012 3952 363018 3964
rect 454494 3952 454500 3964
rect 454552 3952 454558 4004
rect 32398 3884 32404 3936
rect 32456 3924 32462 3936
rect 263962 3924 263968 3936
rect 32456 3896 263968 3924
rect 32456 3884 32462 3896
rect 263962 3884 263968 3896
rect 264020 3884 264026 3936
rect 309042 3884 309048 3936
rect 309100 3924 309106 3936
rect 328454 3924 328460 3936
rect 309100 3896 328460 3924
rect 309100 3884 309106 3896
rect 328454 3884 328460 3896
rect 328512 3884 328518 3936
rect 364334 3884 364340 3936
rect 364392 3924 364398 3936
rect 461578 3924 461584 3936
rect 364392 3896 461584 3924
rect 364392 3884 364398 3896
rect 461578 3884 461584 3896
rect 461636 3884 461642 3936
rect 28902 3816 28908 3868
rect 28960 3856 28966 3868
rect 263686 3856 263692 3868
rect 28960 3828 263692 3856
rect 28960 3816 28966 3828
rect 263686 3816 263692 3828
rect 263744 3816 263750 3868
rect 305546 3816 305552 3868
rect 305604 3856 305610 3868
rect 327166 3856 327172 3868
rect 305604 3828 327172 3856
rect 305604 3816 305610 3828
rect 327166 3816 327172 3828
rect 327224 3816 327230 3868
rect 364426 3816 364432 3868
rect 364484 3856 364490 3868
rect 465166 3856 465172 3868
rect 364484 3828 465172 3856
rect 364484 3816 364490 3828
rect 465166 3816 465172 3828
rect 465224 3816 465230 3868
rect 574738 3816 574744 3868
rect 574796 3856 574802 3868
rect 577406 3856 577412 3868
rect 574796 3828 577412 3856
rect 574796 3816 574802 3828
rect 577406 3816 577412 3828
rect 577464 3816 577470 3868
rect 25314 3748 25320 3800
rect 25372 3788 25378 3800
rect 262306 3788 262312 3800
rect 25372 3760 262312 3788
rect 25372 3748 25378 3760
rect 262306 3748 262312 3760
rect 262364 3748 262370 3800
rect 301958 3748 301964 3800
rect 302016 3788 302022 3800
rect 327074 3788 327080 3800
rect 302016 3760 327080 3788
rect 302016 3748 302022 3760
rect 327074 3748 327080 3760
rect 327132 3748 327138 3800
rect 327994 3748 328000 3800
rect 328052 3788 328058 3800
rect 332686 3788 332692 3800
rect 328052 3760 332692 3788
rect 328052 3748 328058 3760
rect 332686 3748 332692 3760
rect 332744 3748 332750 3800
rect 335446 3748 335452 3800
rect 335504 3788 335510 3800
rect 340966 3788 340972 3800
rect 335504 3760 340972 3788
rect 335504 3748 335510 3760
rect 340966 3748 340972 3760
rect 341024 3748 341030 3800
rect 365714 3748 365720 3800
rect 365772 3788 365778 3800
rect 468662 3788 468668 3800
rect 365772 3760 468668 3788
rect 365772 3748 365778 3760
rect 468662 3748 468668 3760
rect 468720 3748 468726 3800
rect 6454 3680 6460 3732
rect 6512 3720 6518 3732
rect 10318 3720 10324 3732
rect 6512 3692 10324 3720
rect 6512 3680 6518 3692
rect 10318 3680 10324 3692
rect 10376 3680 10382 3732
rect 13538 3680 13544 3732
rect 13596 3720 13602 3732
rect 22738 3720 22744 3732
rect 13596 3692 22744 3720
rect 13596 3680 13602 3692
rect 22738 3680 22744 3692
rect 22796 3680 22802 3732
rect 24210 3680 24216 3732
rect 24268 3720 24274 3732
rect 258074 3720 258080 3732
rect 24268 3692 258080 3720
rect 24268 3680 24274 3692
rect 258074 3680 258080 3692
rect 258132 3680 258138 3732
rect 261202 3720 261208 3732
rect 258276 3692 261208 3720
rect 20622 3612 20628 3664
rect 20680 3652 20686 3664
rect 258276 3652 258304 3692
rect 261202 3680 261208 3692
rect 261260 3680 261266 3732
rect 298462 3680 298468 3732
rect 298520 3720 298526 3732
rect 325970 3720 325976 3732
rect 298520 3692 325976 3720
rect 298520 3680 298526 3692
rect 325970 3680 325976 3692
rect 326028 3680 326034 3732
rect 331582 3680 331588 3732
rect 331640 3720 331646 3732
rect 334066 3720 334072 3732
rect 331640 3692 334072 3720
rect 331640 3680 331646 3692
rect 334066 3680 334072 3692
rect 334124 3680 334130 3732
rect 335722 3680 335728 3732
rect 335780 3720 335786 3732
rect 339862 3720 339868 3732
rect 335780 3692 339868 3720
rect 335780 3680 335786 3692
rect 339862 3680 339868 3692
rect 339920 3680 339926 3732
rect 367094 3680 367100 3732
rect 367152 3720 367158 3732
rect 472250 3720 472256 3732
rect 367152 3692 472256 3720
rect 367152 3680 367158 3692
rect 472250 3680 472256 3692
rect 472308 3680 472314 3732
rect 260926 3652 260932 3664
rect 20680 3624 258304 3652
rect 258368 3624 260932 3652
rect 20680 3612 20686 3624
rect 8754 3544 8760 3596
rect 8812 3584 8818 3596
rect 18598 3584 18604 3596
rect 8812 3556 18604 3584
rect 8812 3544 8818 3556
rect 18598 3544 18604 3556
rect 18656 3544 18662 3596
rect 19426 3544 19432 3596
rect 19484 3584 19490 3596
rect 258368 3584 258396 3624
rect 260926 3612 260932 3624
rect 260984 3612 260990 3664
rect 294874 3612 294880 3664
rect 294932 3652 294938 3664
rect 325786 3652 325792 3664
rect 294932 3624 325792 3652
rect 294932 3612 294938 3624
rect 325786 3612 325792 3624
rect 325844 3612 325850 3664
rect 332686 3612 332692 3664
rect 332744 3652 332750 3664
rect 334158 3652 334164 3664
rect 332744 3624 334164 3652
rect 332744 3612 332750 3624
rect 334158 3612 334164 3624
rect 334216 3612 334222 3664
rect 335630 3612 335636 3664
rect 335688 3652 335694 3664
rect 338666 3652 338672 3664
rect 335688 3624 338672 3652
rect 335688 3612 335694 3624
rect 338666 3612 338672 3624
rect 338724 3612 338730 3664
rect 367186 3612 367192 3664
rect 367244 3652 367250 3664
rect 475746 3652 475752 3664
rect 367244 3624 475752 3652
rect 367244 3612 367250 3624
rect 475746 3612 475752 3624
rect 475804 3612 475810 3664
rect 19484 3556 258396 3584
rect 19484 3544 19490 3556
rect 258442 3544 258448 3596
rect 258500 3584 258506 3596
rect 266722 3584 266728 3596
rect 258500 3556 266728 3584
rect 258500 3544 258506 3556
rect 266722 3544 266728 3556
rect 266780 3544 266786 3596
rect 285674 3544 285680 3596
rect 285732 3584 285738 3596
rect 286042 3584 286048 3596
rect 285732 3556 286048 3584
rect 285732 3544 285738 3556
rect 286042 3544 286048 3556
rect 286100 3544 286106 3596
rect 291378 3544 291384 3596
rect 291436 3584 291442 3596
rect 291436 3556 316034 3584
rect 291436 3544 291442 3556
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 13078 3516 13084 3528
rect 7708 3488 13084 3516
rect 7708 3476 7714 3488
rect 13078 3476 13084 3488
rect 13136 3476 13142 3528
rect 15930 3476 15936 3528
rect 15988 3516 15994 3528
rect 259362 3516 259368 3528
rect 15988 3488 259368 3516
rect 15988 3476 15994 3488
rect 259362 3476 259368 3488
rect 259420 3476 259426 3528
rect 316006 3516 316034 3556
rect 323302 3544 323308 3596
rect 323360 3584 323366 3596
rect 331306 3584 331312 3596
rect 323360 3556 331312 3584
rect 323360 3544 323366 3556
rect 331306 3544 331312 3556
rect 331364 3544 331370 3596
rect 333974 3544 333980 3596
rect 334032 3584 334038 3596
rect 334710 3584 334716 3596
rect 334032 3556 334716 3584
rect 334032 3544 334038 3556
rect 334710 3544 334716 3556
rect 334768 3544 334774 3596
rect 335538 3544 335544 3596
rect 335596 3584 335602 3596
rect 337470 3584 337476 3596
rect 335596 3556 337476 3584
rect 335596 3544 335602 3556
rect 337470 3544 337476 3556
rect 337528 3544 337534 3596
rect 356146 3544 356152 3596
rect 356204 3584 356210 3596
rect 356204 3556 356284 3584
rect 356204 3544 356210 3556
rect 324590 3516 324596 3528
rect 316006 3488 324596 3516
rect 324590 3476 324596 3488
rect 324648 3476 324654 3528
rect 326798 3476 326804 3528
rect 326856 3516 326862 3528
rect 332870 3516 332876 3528
rect 326856 3488 332876 3516
rect 326856 3476 326862 3488
rect 332870 3476 332876 3488
rect 332928 3476 332934 3528
rect 338114 3476 338120 3528
rect 338172 3516 338178 3528
rect 348050 3516 348056 3528
rect 338172 3488 348056 3516
rect 338172 3476 338178 3488
rect 348050 3476 348056 3488
rect 348108 3476 348114 3528
rect 349246 3476 349252 3528
rect 349304 3516 349310 3528
rect 350442 3516 350448 3528
rect 349304 3488 350448 3516
rect 349304 3476 349310 3488
rect 350442 3476 350448 3488
rect 350500 3476 350506 3528
rect 1670 3408 1676 3460
rect 1728 3448 1734 3460
rect 7558 3448 7564 3460
rect 1728 3420 7564 3448
rect 1728 3408 1734 3420
rect 7558 3408 7564 3420
rect 7616 3408 7622 3460
rect 11146 3408 11152 3460
rect 11204 3448 11210 3460
rect 259822 3448 259828 3460
rect 11204 3420 259828 3448
rect 11204 3408 11210 3420
rect 259822 3408 259828 3420
rect 259880 3408 259886 3460
rect 284294 3408 284300 3460
rect 284352 3448 284358 3460
rect 323026 3448 323032 3460
rect 284352 3420 323032 3448
rect 284352 3408 284358 3420
rect 323026 3408 323032 3420
rect 323084 3408 323090 3460
rect 325602 3408 325608 3460
rect 325660 3448 325666 3460
rect 332594 3448 332600 3460
rect 325660 3420 332600 3448
rect 325660 3408 325666 3420
rect 332594 3408 332600 3420
rect 332652 3408 332658 3460
rect 338206 3408 338212 3460
rect 338264 3448 338270 3460
rect 351638 3448 351644 3460
rect 338264 3420 351644 3448
rect 338264 3408 338270 3420
rect 351638 3408 351644 3420
rect 351696 3408 351702 3460
rect 38378 3340 38384 3392
rect 38436 3380 38442 3392
rect 39298 3380 39304 3392
rect 38436 3352 39304 3380
rect 38436 3340 38442 3352
rect 39298 3340 39304 3352
rect 39356 3340 39362 3392
rect 46658 3340 46664 3392
rect 46716 3380 46722 3392
rect 268102 3380 268108 3392
rect 46716 3352 268108 3380
rect 46716 3340 46722 3352
rect 268102 3340 268108 3352
rect 268160 3340 268166 3392
rect 322106 3340 322112 3392
rect 322164 3380 322170 3392
rect 331490 3380 331496 3392
rect 322164 3352 331496 3380
rect 322164 3340 322170 3352
rect 331490 3340 331496 3352
rect 331548 3340 331554 3392
rect 60734 3272 60740 3324
rect 60792 3312 60798 3324
rect 61654 3312 61660 3324
rect 60792 3284 61660 3312
rect 60792 3272 60798 3284
rect 61654 3272 61660 3284
rect 61712 3272 61718 3324
rect 85574 3272 85580 3324
rect 85632 3312 85638 3324
rect 86494 3312 86500 3324
rect 85632 3284 86500 3312
rect 85632 3272 85638 3284
rect 86494 3272 86500 3284
rect 86552 3272 86558 3324
rect 121086 3272 121092 3324
rect 121144 3312 121150 3324
rect 284662 3312 284668 3324
rect 121144 3284 284668 3312
rect 121144 3272 121150 3284
rect 284662 3272 284668 3284
rect 284720 3272 284726 3324
rect 287790 3272 287796 3324
rect 287848 3312 287854 3324
rect 323210 3312 323216 3324
rect 287848 3284 323216 3312
rect 287848 3272 287854 3284
rect 323210 3272 323216 3284
rect 323268 3272 323274 3324
rect 356256 3312 356284 3556
rect 382458 3544 382464 3596
rect 382516 3584 382522 3596
rect 383562 3584 383568 3596
rect 382516 3556 383568 3584
rect 382516 3544 382522 3556
rect 383562 3544 383568 3556
rect 383620 3544 383626 3596
rect 392118 3544 392124 3596
rect 392176 3584 392182 3596
rect 580994 3584 581000 3596
rect 392176 3556 581000 3584
rect 392176 3544 392182 3556
rect 580994 3544 581000 3556
rect 581052 3544 581058 3596
rect 368474 3476 368480 3528
rect 368532 3516 368538 3528
rect 479334 3516 479340 3528
rect 368532 3488 479340 3516
rect 368532 3476 368538 3488
rect 479334 3476 479340 3488
rect 479392 3476 479398 3528
rect 489914 3476 489920 3528
rect 489972 3516 489978 3528
rect 490742 3516 490748 3528
rect 489972 3488 490748 3516
rect 489972 3476 489978 3488
rect 490742 3476 490748 3488
rect 490800 3476 490806 3528
rect 506474 3476 506480 3528
rect 506532 3516 506538 3528
rect 507302 3516 507308 3528
rect 506532 3488 507308 3516
rect 506532 3476 506538 3488
rect 507302 3476 507308 3488
rect 507360 3476 507366 3528
rect 539594 3476 539600 3528
rect 539652 3516 539658 3528
rect 540422 3516 540428 3528
rect 539652 3488 540428 3516
rect 539652 3476 539658 3488
rect 540422 3476 540428 3488
rect 540480 3476 540486 3528
rect 564434 3476 564440 3528
rect 564492 3516 564498 3528
rect 565262 3516 565268 3528
rect 564492 3488 565268 3516
rect 564492 3476 564498 3488
rect 565262 3476 565268 3488
rect 565320 3476 565326 3528
rect 567838 3476 567844 3528
rect 567896 3516 567902 3528
rect 569126 3516 569132 3528
rect 567896 3488 569132 3516
rect 567896 3476 567902 3488
rect 569126 3476 569132 3488
rect 569184 3476 569190 3528
rect 570598 3476 570604 3528
rect 570656 3516 570662 3528
rect 571518 3516 571524 3528
rect 570656 3488 571524 3516
rect 570656 3476 570662 3488
rect 571518 3476 571524 3488
rect 571576 3476 571582 3528
rect 571978 3476 571984 3528
rect 572036 3516 572042 3528
rect 572714 3516 572720 3528
rect 572036 3488 572720 3516
rect 572036 3476 572042 3488
rect 572714 3476 572720 3488
rect 572772 3476 572778 3528
rect 374086 3408 374092 3460
rect 374144 3448 374150 3460
rect 375282 3448 375288 3460
rect 374144 3420 375288 3448
rect 374144 3408 374150 3420
rect 375282 3408 375288 3420
rect 375340 3408 375346 3460
rect 390554 3408 390560 3460
rect 390612 3448 390618 3460
rect 391842 3448 391848 3460
rect 390612 3420 391848 3448
rect 390612 3408 390618 3420
rect 391842 3408 391848 3420
rect 391900 3408 391906 3460
rect 391934 3408 391940 3460
rect 391992 3448 391998 3460
rect 582190 3448 582196 3460
rect 391992 3420 582196 3448
rect 391992 3408 391998 3420
rect 582190 3408 582196 3420
rect 582248 3408 582254 3460
rect 357434 3340 357440 3392
rect 357492 3380 357498 3392
rect 433242 3380 433248 3392
rect 357492 3352 433248 3380
rect 357492 3340 357498 3352
rect 433242 3340 433248 3352
rect 433300 3340 433306 3392
rect 440326 3340 440332 3392
rect 440384 3380 440390 3392
rect 441522 3380 441528 3392
rect 440384 3352 441528 3380
rect 440384 3340 440390 3352
rect 441522 3340 441528 3352
rect 441580 3340 441586 3392
rect 448606 3340 448612 3392
rect 448664 3380 448670 3392
rect 449802 3380 449808 3392
rect 448664 3352 449808 3380
rect 448664 3340 448670 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 572070 3340 572076 3392
rect 572128 3380 572134 3392
rect 573910 3380 573916 3392
rect 572128 3352 573916 3380
rect 572128 3340 572134 3352
rect 573910 3340 573916 3352
rect 573968 3340 573974 3392
rect 356256 3284 423536 3312
rect 124674 3204 124680 3256
rect 124732 3244 124738 3256
rect 285674 3244 285680 3256
rect 124732 3216 285680 3244
rect 124732 3204 124738 3216
rect 285674 3204 285680 3216
rect 285732 3204 285738 3256
rect 329190 3204 329196 3256
rect 329248 3244 329254 3256
rect 332778 3244 332784 3256
rect 329248 3216 332784 3244
rect 329248 3204 329254 3216
rect 332778 3204 332784 3216
rect 332836 3204 332842 3256
rect 356422 3204 356428 3256
rect 356480 3244 356486 3256
rect 356480 3216 412634 3244
rect 356480 3204 356486 3216
rect 258074 3136 258080 3188
rect 258132 3176 258138 3188
rect 262582 3176 262588 3188
rect 258132 3148 262588 3176
rect 258132 3136 258138 3148
rect 262582 3136 262588 3148
rect 262640 3136 262646 3188
rect 330386 3136 330392 3188
rect 330444 3176 330450 3188
rect 334342 3176 334348 3188
rect 330444 3148 334348 3176
rect 330444 3136 330450 3148
rect 334342 3136 334348 3148
rect 334400 3136 334406 3188
rect 398926 3136 398932 3188
rect 398984 3176 398990 3188
rect 400122 3176 400128 3188
rect 398984 3148 400128 3176
rect 398984 3136 398990 3148
rect 400122 3136 400128 3148
rect 400180 3136 400186 3188
rect 407206 3136 407212 3188
rect 407264 3176 407270 3188
rect 408402 3176 408408 3188
rect 407264 3148 408408 3176
rect 407264 3136 407270 3148
rect 408402 3136 408408 3148
rect 408460 3136 408466 3188
rect 566 3068 572 3120
rect 624 3108 630 3120
rect 4798 3108 4804 3120
rect 624 3080 4804 3108
rect 624 3068 630 3080
rect 4798 3068 4804 3080
rect 4856 3068 4862 3120
rect 23014 3068 23020 3120
rect 23072 3108 23078 3120
rect 25498 3108 25504 3120
rect 23072 3080 25504 3108
rect 23072 3068 23078 3080
rect 25498 3068 25504 3080
rect 25556 3068 25562 3120
rect 412606 3108 412634 3216
rect 415394 3204 415400 3256
rect 415452 3244 415458 3256
rect 416682 3244 416688 3256
rect 415452 3216 416688 3244
rect 415452 3204 415458 3216
rect 416682 3204 416688 3216
rect 416740 3204 416746 3256
rect 423508 3176 423536 3284
rect 423674 3272 423680 3324
rect 423732 3312 423738 3324
rect 424962 3312 424968 3324
rect 423732 3284 424968 3312
rect 423732 3272 423738 3284
rect 424962 3272 424968 3284
rect 425020 3272 425026 3324
rect 429654 3176 429660 3188
rect 423508 3148 429660 3176
rect 429654 3136 429660 3148
rect 429712 3136 429718 3188
rect 426158 3108 426164 3120
rect 412606 3080 426164 3108
rect 426158 3068 426164 3080
rect 426216 3068 426222 3120
rect 12342 3000 12348 3052
rect 12400 3040 12406 3052
rect 14458 3040 14464 3052
rect 12400 3012 14464 3040
rect 12400 3000 12406 3012
rect 14458 3000 14464 3012
rect 14516 3000 14522 3052
rect 336826 3000 336832 3052
rect 336884 3040 336890 3052
rect 344554 3040 344560 3052
rect 336884 3012 344560 3040
rect 336884 3000 336890 3012
rect 344554 3000 344560 3012
rect 344612 3000 344618 3052
rect 336734 2932 336740 2984
rect 336792 2972 336798 2984
rect 343358 2972 343364 2984
rect 336792 2944 343364 2972
rect 336792 2932 336798 2944
rect 343358 2932 343364 2944
rect 343416 2932 343422 2984
rect 456794 1640 456800 1692
rect 456852 1680 456858 1692
rect 458082 1680 458088 1692
rect 456852 1652 458088 1680
rect 456852 1640 456858 1652
rect 458082 1640 458088 1652
rect 458140 1640 458146 1692
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 322940 700748 322992 700800
rect 348792 700748 348844 700800
rect 283840 700680 283892 700732
rect 328460 700680 328512 700732
rect 318800 700612 318852 700664
rect 413652 700612 413704 700664
rect 218980 700544 219032 700596
rect 332600 700544 332652 700596
rect 154120 700476 154172 700528
rect 338120 700476 338172 700528
rect 89168 700408 89220 700460
rect 342260 700408 342312 700460
rect 24308 700340 24360 700392
rect 346400 700340 346452 700392
rect 8116 700272 8168 700324
rect 345020 700272 345072 700324
rect 413284 700272 413336 700324
rect 559656 700272 559708 700324
rect 300124 700000 300176 700052
rect 301504 700000 301556 700052
rect 105452 699660 105504 699712
rect 106924 699660 106976 699712
rect 428464 699660 428516 699712
rect 429844 699660 429896 699712
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 303620 696940 303672 696992
rect 580172 696940 580224 696992
rect 305000 683136 305052 683188
rect 580172 683136 580224 683188
rect 302240 670760 302292 670812
rect 580172 670760 580224 670812
rect 3516 670692 3568 670744
rect 351920 670692 351972 670744
rect 3516 656888 3568 656940
rect 350540 656888 350592 656940
rect 298100 643084 298152 643136
rect 580172 643084 580224 643136
rect 299480 630640 299532 630692
rect 580172 630640 580224 630692
rect 3332 618264 3384 618316
rect 356060 618264 356112 618316
rect 296720 616836 296772 616888
rect 580172 616836 580224 616888
rect 3332 605820 3384 605872
rect 354680 605820 354732 605872
rect 293960 590656 294012 590708
rect 579804 590656 579856 590708
rect 295340 576852 295392 576904
rect 580172 576852 580224 576904
rect 3056 565836 3108 565888
rect 361580 565836 361632 565888
rect 292580 563048 292632 563100
rect 579804 563048 579856 563100
rect 3332 553392 3384 553444
rect 358820 553392 358872 553444
rect 288440 536800 288492 536852
rect 580172 536800 580224 536852
rect 291200 524424 291252 524476
rect 580172 524424 580224 524476
rect 3332 514768 3384 514820
rect 365720 514768 365772 514820
rect 287060 510620 287112 510672
rect 580172 510620 580224 510672
rect 320180 502936 320232 502988
rect 364340 502936 364392 502988
rect 3240 500964 3292 501016
rect 364340 500964 364392 501016
rect 284300 484372 284352 484424
rect 580172 484372 580224 484424
rect 40040 473968 40092 474020
rect 344100 473968 344152 474020
rect 311256 472608 311308 472660
rect 494060 472608 494112 472660
rect 286232 470568 286284 470620
rect 579988 470568 580040 470620
rect 106924 469820 106976 469872
rect 339500 469820 339552 469872
rect 169760 468460 169812 468512
rect 334716 468460 334768 468512
rect 234620 467100 234672 467152
rect 330024 467100 330076 467152
rect 301504 465672 301556 465724
rect 325700 465672 325752 465724
rect 316040 464312 316092 464364
rect 428464 464312 428516 464364
rect 277216 464040 277268 464092
rect 435364 464040 435416 464092
rect 215944 463972 215996 464024
rect 380072 463972 380124 464024
rect 220084 463904 220136 463956
rect 387892 463904 387944 463956
rect 217324 463836 217376 463888
rect 392584 463836 392636 463888
rect 280712 463768 280764 463820
rect 457444 463768 457496 463820
rect 13084 463700 13136 463752
rect 378508 463700 378560 463752
rect 235356 462816 235408 462868
rect 375472 462816 375524 462868
rect 264888 462748 264940 462800
rect 422944 462748 422996 462800
rect 221464 462680 221516 462732
rect 383292 462680 383344 462732
rect 260380 462612 260432 462664
rect 421564 462612 421616 462664
rect 279148 462544 279200 462596
rect 454684 462544 454736 462596
rect 247868 462476 247920 462528
rect 427084 462476 427136 462528
rect 242808 462408 242860 462460
rect 424324 462408 424376 462460
rect 3516 462340 3568 462392
rect 370780 462340 370832 462392
rect 307300 461592 307352 461644
rect 413284 461592 413336 461644
rect 236736 461388 236788 461440
rect 374000 461388 374052 461440
rect 229744 461320 229796 461372
rect 396080 461320 396132 461372
rect 250904 461252 250956 461304
rect 417424 461252 417476 461304
rect 257252 461184 257304 461236
rect 428464 461184 428516 461236
rect 228364 461116 228416 461168
rect 400496 461116 400548 461168
rect 224224 461048 224276 461100
rect 409880 461048 409932 461100
rect 269764 460980 269816 461032
rect 567936 460980 567988 461032
rect 18696 460912 18748 460964
rect 391112 460912 391164 460964
rect 201500 460844 201552 460896
rect 331680 460844 331732 460896
rect 313188 460776 313240 460828
rect 462320 460776 462372 460828
rect 315120 460708 315172 460760
rect 477500 460708 477552 460760
rect 136640 460640 136692 460692
rect 336372 460640 336424 460692
rect 308864 460572 308916 460624
rect 527180 460572 527232 460624
rect 310428 460504 310480 460556
rect 542360 460504 542412 460556
rect 71780 460436 71832 460488
rect 341064 460436 341116 460488
rect 3608 460368 3660 460420
rect 353576 460368 353628 460420
rect 3700 460300 3752 460352
rect 358268 460300 358320 460352
rect 3792 460232 3844 460284
rect 362960 460232 363012 460284
rect 3884 460164 3936 460216
rect 367652 460164 367704 460216
rect 318248 460096 318300 460148
rect 397460 460096 397512 460148
rect 266360 460028 266412 460080
rect 327080 460028 327132 460080
rect 322848 459960 322900 460012
rect 331220 459960 331272 460012
rect 282276 459552 282328 459604
rect 308496 459552 308548 459604
rect 353300 459552 353352 459604
rect 369216 459552 369268 459604
rect 235264 458872 235316 458924
rect 377036 458872 377088 458924
rect 308496 458804 308548 458856
rect 580356 458804 580408 458856
rect 274456 458736 274508 458788
rect 416044 458736 416096 458788
rect 233976 458668 234028 458720
rect 381728 458668 381780 458720
rect 232504 458600 232556 458652
rect 386420 458600 386472 458652
rect 255688 458532 255740 458584
rect 418804 458532 418856 458584
rect 266268 458464 266320 458516
rect 431224 458464 431276 458516
rect 246304 458396 246356 458448
rect 414664 458396 414716 458448
rect 225604 458328 225656 458380
rect 405188 458328 405240 458380
rect 241428 458260 241480 458312
rect 580264 458260 580316 458312
rect 3424 458192 3476 458244
rect 372666 458192 372718 458244
rect 238024 457512 238076 457564
rect 239404 457512 239456 457564
rect 3516 457444 3568 457496
rect 275928 457444 275980 457496
rect 283656 457444 283708 457496
rect 353300 457444 353352 457496
rect 412088 457444 412140 457496
rect 414112 457444 414164 457496
rect 432604 456832 432656 456884
rect 580172 456764 580224 456816
rect 457444 431876 457496 431928
rect 579620 431876 579672 431928
rect 3424 411204 3476 411256
rect 235356 411204 235408 411256
rect 454684 405628 454736 405680
rect 579620 405628 579672 405680
rect 3240 398760 3292 398812
rect 235908 398760 235960 398812
rect 432604 379448 432656 379500
rect 580172 379448 580224 379500
rect 3240 372512 3292 372564
rect 235264 372512 235316 372564
rect 435364 365644 435416 365696
rect 580172 365644 580224 365696
rect 3332 358708 3384 358760
rect 215944 358708 215996 358760
rect 416044 353200 416096 353252
rect 580172 353200 580224 353252
rect 3148 346332 3200 346384
rect 13084 346332 13136 346384
rect 256056 336676 256108 336728
rect 257804 336676 257856 336728
rect 264244 336676 264296 336728
rect 266360 336676 266412 336728
rect 271144 336676 271196 336728
rect 273260 336676 273312 336728
rect 273904 336676 273956 336728
rect 275008 336676 275060 336728
rect 278872 336676 278924 336728
rect 279148 336676 279200 336728
rect 279424 336676 279476 336728
rect 280436 336676 280488 336728
rect 284484 336676 284536 336728
rect 284852 336676 284904 336728
rect 287704 336676 287756 336728
rect 288992 336676 289044 336728
rect 289176 336676 289228 336728
rect 290372 336676 290424 336728
rect 293224 336676 293276 336728
rect 294236 336676 294288 336728
rect 296812 336676 296864 336728
rect 297548 336676 297600 336728
rect 298744 336676 298796 336728
rect 300032 336676 300084 336728
rect 300860 336676 300912 336728
rect 301136 336676 301188 336728
rect 302240 336676 302292 336728
rect 302516 336676 302568 336728
rect 303620 336676 303672 336728
rect 303988 336676 304040 336728
rect 309876 336676 309928 336728
rect 312728 336676 312780 336728
rect 318892 336676 318944 336728
rect 319076 336676 319128 336728
rect 327724 336676 327776 336728
rect 331220 336676 331272 336728
rect 334072 336676 334124 336728
rect 334348 336676 334400 336728
rect 336740 336676 336792 336728
rect 337108 336676 337160 336728
rect 348608 336676 348660 336728
rect 349804 336676 349856 336728
rect 353484 336676 353536 336728
rect 353668 336676 353720 336728
rect 356244 336676 356296 336728
rect 356428 336676 356480 336728
rect 372712 336676 372764 336728
rect 372988 336676 373040 336728
rect 376208 336676 376260 336728
rect 377404 336676 377456 336728
rect 378324 336676 378376 336728
rect 378508 336676 378560 336728
rect 386604 336676 386656 336728
rect 386788 336676 386840 336728
rect 256148 336608 256200 336660
rect 260840 336608 260892 336660
rect 268384 336608 268436 336660
rect 272156 336608 272208 336660
rect 303528 336608 303580 336660
rect 311900 336608 311952 336660
rect 318064 336608 318116 336660
rect 320456 336608 320508 336660
rect 257344 336540 257396 336592
rect 268844 336540 268896 336592
rect 305736 336540 305788 336592
rect 316040 336540 316092 336592
rect 316684 336540 316736 336592
rect 322112 336540 322164 336592
rect 348700 336540 348752 336592
rect 370504 336540 370556 336592
rect 377496 336540 377548 336592
rect 399484 336540 399536 336592
rect 233884 336472 233936 336524
rect 264704 336472 264756 336524
rect 307024 336472 307076 336524
rect 322940 336472 322992 336524
rect 323584 336472 323636 336524
rect 324596 336472 324648 336524
rect 344284 336472 344336 336524
rect 359556 336472 359608 336524
rect 370780 336472 370832 336524
rect 395344 336472 395396 336524
rect 255964 336404 256016 336456
rect 296168 336404 296220 336456
rect 301504 336404 301556 336456
rect 317696 336404 317748 336456
rect 342076 336404 342128 336456
rect 363604 336404 363656 336456
rect 369952 336404 370004 336456
rect 396724 336404 396776 336456
rect 243544 336336 243596 336388
rect 287888 336336 287940 336388
rect 305644 336336 305696 336388
rect 323492 336336 323544 336388
rect 346768 336336 346820 336388
rect 378784 336336 378836 336388
rect 382372 336336 382424 336388
rect 407764 336336 407816 336388
rect 242164 336268 242216 336320
rect 296444 336268 296496 336320
rect 304264 336268 304316 336320
rect 322664 336268 322716 336320
rect 340052 336268 340104 336320
rect 341524 336268 341576 336320
rect 345112 336268 345164 336320
rect 371884 336268 371936 336320
rect 374276 336268 374328 336320
rect 410524 336268 410576 336320
rect 247684 336200 247736 336252
rect 307760 336200 307812 336252
rect 309784 336200 309836 336252
rect 320180 336200 320232 336252
rect 322204 336200 322256 336252
rect 330944 336200 330996 336252
rect 340144 336200 340196 336252
rect 356060 336200 356112 336252
rect 358912 336200 358964 336252
rect 436100 336200 436152 336252
rect 117320 336132 117372 336184
rect 284300 336132 284352 336184
rect 297548 336132 297600 336184
rect 298652 336132 298704 336184
rect 300124 336132 300176 336184
rect 321836 336132 321888 336184
rect 360568 336132 360620 336184
rect 443000 336132 443052 336184
rect 110420 336064 110472 336116
rect 282644 336064 282696 336116
rect 295984 336064 296036 336116
rect 319352 336064 319404 336116
rect 320824 336064 320876 336116
rect 330116 336064 330168 336116
rect 342352 336064 342404 336116
rect 360844 336064 360896 336116
rect 362224 336064 362276 336116
rect 449900 336064 449952 336116
rect 10324 335996 10376 336048
rect 269764 335996 269816 336048
rect 271052 335996 271104 336048
rect 285680 335996 285732 336048
rect 294512 335996 294564 336048
rect 297180 335996 297232 336048
rect 324320 335996 324372 336048
rect 341248 335996 341300 336048
rect 359464 335996 359516 336048
rect 363880 335996 363932 336048
rect 456800 335996 456852 336048
rect 258356 335928 258408 335980
rect 284300 335928 284352 335980
rect 286232 335928 286284 335980
rect 293316 335928 293368 335980
rect 293960 335928 294012 335980
rect 356704 335860 356756 335912
rect 360568 335860 360620 335912
rect 365812 335860 365864 335912
rect 369124 335860 369176 335912
rect 271236 335792 271288 335844
rect 272984 335792 273036 335844
rect 343732 335792 343784 335844
rect 345664 335792 345716 335844
rect 357532 335724 357584 335776
rect 360936 335724 360988 335776
rect 261484 335656 261536 335708
rect 263048 335656 263100 335708
rect 275284 335656 275336 335708
rect 276296 335656 276348 335708
rect 287796 335656 287848 335708
rect 288716 335656 288768 335708
rect 291844 335656 291896 335708
rect 293132 335656 293184 335708
rect 315304 335656 315356 335708
rect 317144 335656 317196 335708
rect 361672 335656 361724 335708
rect 363696 335656 363748 335708
rect 297456 335588 297508 335640
rect 298100 335588 298152 335640
rect 289084 335520 289136 335572
rect 289820 335520 289872 335572
rect 296168 335452 296220 335504
rect 298376 335452 298428 335504
rect 311164 335452 311216 335504
rect 317972 335452 318024 335504
rect 296076 335384 296128 335436
rect 297272 335384 297324 335436
rect 323676 335384 323728 335436
rect 326804 335384 326856 335436
rect 392032 335384 392084 335436
rect 393964 335384 394016 335436
rect 257436 335316 257488 335368
rect 259184 335316 259236 335368
rect 286324 335316 286376 335368
rect 287612 335316 287664 335368
rect 296260 335316 296312 335368
rect 296996 335316 297048 335368
rect 302884 335316 302936 335368
rect 306656 335316 306708 335368
rect 313924 335316 313976 335368
rect 316868 335316 316920 335368
rect 324964 335316 325016 335368
rect 325976 335316 326028 335368
rect 283196 335248 283248 335300
rect 283380 335248 283432 335300
rect 332876 335248 332928 335300
rect 333060 335248 333112 335300
rect 234620 334772 234672 334824
rect 303528 334772 303580 334824
rect 205640 334704 205692 334756
rect 305000 334704 305052 334756
rect 359372 334704 359424 334756
rect 438860 334704 438912 334756
rect 160100 334636 160152 334688
rect 285680 334636 285732 334688
rect 369216 334636 369268 334688
rect 480260 334636 480312 334688
rect 14464 334568 14516 334620
rect 259828 334568 259880 334620
rect 380808 334568 380860 334620
rect 529940 334568 529992 334620
rect 248420 333412 248472 333464
rect 314936 333412 314988 333464
rect 220820 333344 220872 333396
rect 308588 333344 308640 333396
rect 360476 333344 360528 333396
rect 441620 333344 441672 333396
rect 125600 333276 125652 333328
rect 284300 333276 284352 333328
rect 13084 333208 13136 333260
rect 258632 333140 258684 333192
rect 372528 333072 372580 333124
rect 494060 333276 494112 333328
rect 384948 333208 385000 333260
rect 547880 333208 547932 333260
rect 242900 331984 242952 332036
rect 313832 331984 313884 332036
rect 349620 331984 349672 332036
rect 396080 331984 396132 332036
rect 207020 331916 207072 331968
rect 305368 331916 305420 331968
rect 371700 331916 371752 331968
rect 489920 331916 489972 331968
rect 98000 331848 98052 331900
rect 279884 331848 279936 331900
rect 384212 331848 384264 331900
rect 543740 331848 543792 331900
rect 377036 331168 377088 331220
rect 377220 331168 377272 331220
rect 327356 330896 327408 330948
rect 292764 330692 292816 330744
rect 292948 330692 293000 330744
rect 253940 330624 253992 330676
rect 316316 330624 316368 330676
rect 334348 330760 334400 330812
rect 352012 330624 352064 330676
rect 407120 330624 407172 330676
rect 213920 330556 213972 330608
rect 306932 330556 306984 330608
rect 327356 330556 327408 330608
rect 334348 330556 334400 330608
rect 373356 330556 373408 330608
rect 498200 330556 498252 330608
rect 103520 330488 103572 330540
rect 273444 330420 273496 330472
rect 274088 330420 274140 330472
rect 274824 330420 274876 330472
rect 275468 330420 275520 330472
rect 277400 330420 277452 330472
rect 278228 330420 278280 330472
rect 278964 330488 279016 330540
rect 279608 330488 279660 330540
rect 281632 330488 281684 330540
rect 282368 330488 282420 330540
rect 282920 330488 282972 330540
rect 283472 330488 283524 330540
rect 284392 330488 284444 330540
rect 285404 330488 285456 330540
rect 285956 330488 286008 330540
rect 286508 330488 286560 330540
rect 287336 330488 287388 330540
rect 288164 330488 288216 330540
rect 288716 330488 288768 330540
rect 289268 330488 289320 330540
rect 291568 330488 291620 330540
rect 292304 330488 292356 330540
rect 292672 330488 292724 330540
rect 293684 330488 293736 330540
rect 296996 330488 297048 330540
rect 297824 330488 297876 330540
rect 298192 330488 298244 330540
rect 298928 330488 298980 330540
rect 301136 330488 301188 330540
rect 301964 330488 302016 330540
rect 313648 330488 313700 330540
rect 314108 330488 314160 330540
rect 317696 330488 317748 330540
rect 318248 330488 318300 330540
rect 321652 330488 321704 330540
rect 322388 330488 322440 330540
rect 323216 330488 323268 330540
rect 324044 330488 324096 330540
rect 324412 330488 324464 330540
rect 325148 330488 325200 330540
rect 327172 330488 327224 330540
rect 328184 330488 328236 330540
rect 328736 330488 328788 330540
rect 329564 330488 329616 330540
rect 331312 330488 331364 330540
rect 332324 330488 332376 330540
rect 332692 330488 332744 330540
rect 333428 330488 333480 330540
rect 334256 330488 334308 330540
rect 334808 330488 334860 330540
rect 335452 330488 335504 330540
rect 336464 330488 336516 330540
rect 336832 330488 336884 330540
rect 337292 330488 337344 330540
rect 338212 330488 338264 330540
rect 338948 330488 339000 330540
rect 339500 330488 339552 330540
rect 340604 330488 340656 330540
rect 360292 330488 360344 330540
rect 361028 330488 361080 330540
rect 361580 330488 361632 330540
rect 362684 330488 362736 330540
rect 363144 330488 363196 330540
rect 364064 330488 364116 330540
rect 364524 330488 364576 330540
rect 365168 330488 365220 330540
rect 365720 330488 365772 330540
rect 366272 330488 366324 330540
rect 368480 330488 368532 330540
rect 368756 330488 368808 330540
rect 389456 330488 389508 330540
rect 390008 330488 390060 330540
rect 390836 330488 390888 330540
rect 391664 330488 391716 330540
rect 391940 330488 391992 330540
rect 392492 330488 392544 330540
rect 281264 330420 281316 330472
rect 283012 330420 283064 330472
rect 284024 330420 284076 330472
rect 285864 330420 285916 330472
rect 286784 330420 286836 330472
rect 288624 330420 288676 330472
rect 289544 330420 289596 330472
rect 292856 330420 292908 330472
rect 293408 330420 293460 330472
rect 298284 330420 298336 330472
rect 299204 330420 299256 330472
rect 313464 330420 313516 330472
rect 314384 330420 314436 330472
rect 315028 330420 315080 330472
rect 315488 330420 315540 330472
rect 317512 330420 317564 330472
rect 318524 330420 318576 330472
rect 324504 330420 324556 330472
rect 325424 330420 325476 330472
rect 327448 330420 327500 330472
rect 327908 330420 327960 330472
rect 328460 330420 328512 330472
rect 329012 330420 329064 330472
rect 332876 330420 332928 330472
rect 333152 330420 333204 330472
rect 333980 330420 334032 330472
rect 335084 330420 335136 330472
rect 336924 330420 336976 330472
rect 337568 330420 337620 330472
rect 338304 330420 338356 330472
rect 339224 330420 339276 330472
rect 360200 330420 360252 330472
rect 361304 330420 361356 330472
rect 364432 330420 364484 330472
rect 365444 330420 365496 330472
rect 365812 330420 365864 330472
rect 366824 330420 366876 330472
rect 368572 330420 368624 330472
rect 369584 330420 369636 330472
rect 392032 330420 392084 330472
rect 392768 330420 392820 330472
rect 273352 330352 273404 330404
rect 274364 330352 274416 330404
rect 274732 330352 274784 330404
rect 275744 330352 275796 330404
rect 283196 330352 283248 330404
rect 283748 330352 283800 330404
rect 299848 330352 299900 330404
rect 300584 330352 300636 330404
rect 390560 330352 390612 330404
rect 571984 330488 572036 330540
rect 299664 330284 299716 330336
rect 300308 330284 300360 330336
rect 332784 330148 332836 330200
rect 333704 330148 333756 330200
rect 277676 329808 277728 329860
rect 277952 329808 278004 329860
rect 323124 329740 323176 329792
rect 323768 329740 323820 329792
rect 389272 329400 389324 329452
rect 390284 329400 390336 329452
rect 277584 329264 277636 329316
rect 278504 329264 278556 329316
rect 360568 329196 360620 329248
rect 426440 329196 426492 329248
rect 224960 329128 225012 329180
rect 309600 329128 309652 329180
rect 375932 329128 375984 329180
rect 507860 329128 507912 329180
rect 149060 329060 149112 329112
rect 291752 329060 291804 329112
rect 384396 329060 384448 329112
rect 545120 329060 545172 329112
rect 364248 328516 364300 328568
rect 364708 328516 364760 328568
rect 311992 328312 312044 328364
rect 313004 328312 313056 328364
rect 367192 328176 367244 328228
rect 367928 328176 367980 328228
rect 320456 328040 320508 328092
rect 321284 328040 321336 328092
rect 339592 328040 339644 328092
rect 340328 328040 340380 328092
rect 361672 327904 361724 327956
rect 362408 327904 362460 327956
rect 189080 327836 189132 327888
rect 300860 327836 300912 327888
rect 161480 327768 161532 327820
rect 294788 327768 294840 327820
rect 363696 327768 363748 327820
rect 448520 327768 448572 327820
rect 85580 327700 85632 327752
rect 277124 327700 277176 327752
rect 314752 327700 314804 327752
rect 315764 327700 315816 327752
rect 376484 327700 376536 327752
rect 512000 327700 512052 327752
rect 291292 327020 291344 327072
rect 292028 327020 292080 327072
rect 319076 326884 319128 326936
rect 319904 326884 319956 326936
rect 269396 326680 269448 326732
rect 269580 326680 269632 326732
rect 363052 326612 363104 326664
rect 363512 326612 363564 326664
rect 263784 326544 263836 326596
rect 264060 326544 264112 326596
rect 269304 326544 269356 326596
rect 269488 326544 269540 326596
rect 320272 326544 320324 326596
rect 321008 326544 321060 326596
rect 201500 326476 201552 326528
rect 303620 326476 303672 326528
rect 382372 326476 382424 326528
rect 383384 326476 383436 326528
rect 385316 326476 385368 326528
rect 385500 326476 385552 326528
rect 182180 326408 182232 326460
rect 299480 326408 299532 326460
rect 302332 326408 302384 326460
rect 303344 326408 303396 326460
rect 303988 326408 304040 326460
rect 304448 326408 304500 326460
rect 305184 326408 305236 326460
rect 306104 326408 306156 326460
rect 309324 326408 309376 326460
rect 310244 326408 310296 326460
rect 345204 326408 345256 326460
rect 346124 326408 346176 326460
rect 346400 326408 346452 326460
rect 347504 326408 347556 326460
rect 347964 326408 348016 326460
rect 348148 326408 348200 326460
rect 350724 326408 350776 326460
rect 351000 326408 351052 326460
rect 353392 326408 353444 326460
rect 354404 326408 354456 326460
rect 354772 326408 354824 326460
rect 355508 326408 355560 326460
rect 357532 326408 357584 326460
rect 358268 326408 358320 326460
rect 358912 326408 358964 326460
rect 359924 326408 359976 326460
rect 364892 326408 364944 326460
rect 462320 326408 462372 326460
rect 53840 326340 53892 326392
rect 256792 326340 256844 326392
rect 257528 326340 257580 326392
rect 258172 326340 258224 326392
rect 258908 326340 258960 326392
rect 259644 326340 259696 326392
rect 260288 326340 260340 326392
rect 261208 326340 261260 326392
rect 261668 326340 261720 326392
rect 262312 326340 262364 326392
rect 262772 326340 262824 326392
rect 264980 326340 265032 326392
rect 265440 326340 265492 326392
rect 266452 326340 266504 326392
rect 267464 326340 267516 326392
rect 267832 326340 267884 326392
rect 268568 326340 268620 326392
rect 269488 326340 269540 326392
rect 269948 326340 270000 326392
rect 270868 326340 270920 326392
rect 271604 326340 271656 326392
rect 302608 326340 302660 326392
rect 303068 326340 303120 326392
rect 303804 326340 303856 326392
rect 304172 326340 304224 326392
rect 305276 326340 305328 326392
rect 305828 326340 305880 326392
rect 306656 326340 306708 326392
rect 307484 326340 307536 326392
rect 307852 326340 307904 326392
rect 308312 326340 308364 326392
rect 309508 326340 309560 326392
rect 309968 326340 310020 326392
rect 340972 326340 341024 326392
rect 341708 326340 341760 326392
rect 342352 326340 342404 326392
rect 343364 326340 343416 326392
rect 343640 326340 343692 326392
rect 344744 326340 344796 326392
rect 345112 326340 345164 326392
rect 345572 326340 345624 326392
rect 346492 326340 346544 326392
rect 347228 326340 347280 326392
rect 347780 326340 347832 326392
rect 348884 326340 348936 326392
rect 349160 326340 349212 326392
rect 350264 326340 350316 326392
rect 350632 326340 350684 326392
rect 351368 326340 351420 326392
rect 351920 326340 351972 326392
rect 353024 326340 353076 326392
rect 353300 326340 353352 326392
rect 353852 326340 353904 326392
rect 354956 326340 355008 326392
rect 355232 326340 355284 326392
rect 356152 326340 356204 326392
rect 357164 326340 357216 326392
rect 357440 326340 357492 326392
rect 357992 326340 358044 326392
rect 358820 326340 358872 326392
rect 359648 326340 359700 326392
rect 369860 326340 369912 326392
rect 370412 326340 370464 326392
rect 371332 326340 371384 326392
rect 372068 326340 372120 326392
rect 372896 326340 372948 326392
rect 373448 326340 373500 326392
rect 374184 326340 374236 326392
rect 374552 326340 374604 326392
rect 375380 326340 375432 326392
rect 376300 326340 376352 326392
rect 378232 326340 378284 326392
rect 378968 326340 379020 326392
rect 379520 326340 379572 326392
rect 380348 326340 380400 326392
rect 381084 326340 381136 326392
rect 381728 326340 381780 326392
rect 382464 326340 382516 326392
rect 383108 326340 383160 326392
rect 383660 326340 383712 326392
rect 384488 326340 384540 326392
rect 385040 326340 385092 326392
rect 385868 326340 385920 326392
rect 386696 326340 386748 326392
rect 387248 326340 387300 326392
rect 388076 326340 388128 326392
rect 388904 326340 388956 326392
rect 259552 326204 259604 326256
rect 260564 326204 260616 326256
rect 260932 326204 260984 326256
rect 261392 326204 261444 326256
rect 262404 326204 262456 326256
rect 263324 326204 263376 326256
rect 263968 326204 264020 326256
rect 264428 326204 264480 326256
rect 265164 326204 265216 326256
rect 265808 326204 265860 326256
rect 267924 326204 267976 326256
rect 268292 326204 268344 326256
rect 269212 326272 269264 326324
rect 270224 326272 270276 326324
rect 270776 326272 270828 326324
rect 271328 326272 271380 326324
rect 303712 326272 303764 326324
rect 304724 326272 304776 326324
rect 345020 326272 345072 326324
rect 345848 326272 345900 326324
rect 357624 326272 357676 326324
rect 358544 326272 358596 326324
rect 369952 326272 370004 326324
rect 370964 326272 371016 326324
rect 372804 326272 372856 326324
rect 373724 326272 373776 326324
rect 374276 326272 374328 326324
rect 375104 326272 375156 326324
rect 378140 326272 378192 326324
rect 379244 326272 379296 326324
rect 380992 326272 381044 326324
rect 382004 326272 382056 326324
rect 382280 326272 382332 326324
rect 382832 326272 382884 326324
rect 385132 326272 385184 326324
rect 386144 326272 386196 326324
rect 386420 326272 386472 326324
rect 386972 326272 387024 326324
rect 269672 326204 269724 326256
rect 310612 326204 310664 326256
rect 310796 326204 310848 326256
rect 310888 326204 310940 326256
rect 311624 326204 311676 326256
rect 350816 326204 350868 326256
rect 351644 326204 351696 326256
rect 376944 326204 376996 326256
rect 377588 326204 377640 326256
rect 379796 326204 379848 326256
rect 525800 326340 525852 326392
rect 265072 326136 265124 326188
rect 266084 326136 266136 326188
rect 289912 326136 289964 326188
rect 290648 326136 290700 326188
rect 376852 326136 376904 326188
rect 377864 326136 377916 326188
rect 328552 325864 328604 325916
rect 329288 325864 329340 325916
rect 368756 325864 368808 325916
rect 369308 325864 369360 325916
rect 396816 325592 396868 325644
rect 579896 325592 579948 325644
rect 266636 325320 266688 325372
rect 267188 325320 267240 325372
rect 309232 325320 309284 325372
rect 309692 325320 309744 325372
rect 231860 325048 231912 325100
rect 311072 325048 311124 325100
rect 349804 325048 349856 325100
rect 390560 325048 390612 325100
rect 164240 324980 164292 325032
rect 295340 324980 295392 325032
rect 352472 324980 352524 325032
rect 408500 324980 408552 325032
rect 46940 324912 46992 324964
rect 268108 324912 268160 324964
rect 377220 324912 377272 324964
rect 513380 324912 513432 324964
rect 386512 324640 386564 324692
rect 387524 324640 387576 324692
rect 261116 324504 261168 324556
rect 261944 324504 261996 324556
rect 343732 324368 343784 324420
rect 344468 324368 344520 324420
rect 387800 324300 387852 324352
rect 388628 324300 388680 324352
rect 310612 324232 310664 324284
rect 311348 324232 311400 324284
rect 380900 324096 380952 324148
rect 381268 324096 381320 324148
rect 238760 323756 238812 323808
rect 309876 323756 309928 323808
rect 171140 323688 171192 323740
rect 296260 323688 296312 323740
rect 306472 323688 306524 323740
rect 307208 323688 307260 323740
rect 353668 323688 353720 323740
rect 412640 323688 412692 323740
rect 155960 323620 156012 323672
rect 292856 323620 292908 323672
rect 374828 323620 374880 323672
rect 505100 323620 505152 323672
rect 25504 323552 25556 323604
rect 262496 323552 262548 323604
rect 342444 323552 342496 323604
rect 343088 323552 343140 323604
rect 359556 323552 359608 323604
rect 374000 323552 374052 323604
rect 380072 323552 380124 323604
rect 527180 323552 527232 323604
rect 387984 323212 388036 323264
rect 388352 323212 388404 323264
rect 356336 323144 356388 323196
rect 356888 323144 356940 323196
rect 354680 322736 354732 322788
rect 355784 322736 355836 322788
rect 242992 322396 243044 322448
rect 313556 322396 313608 322448
rect 175280 322328 175332 322380
rect 296996 322328 297048 322380
rect 349252 322328 349304 322380
rect 394700 322328 394752 322380
rect 142160 322260 142212 322312
rect 290004 322260 290056 322312
rect 366548 322260 366600 322312
rect 469220 322260 469272 322312
rect 34520 322192 34572 322244
rect 265348 322192 265400 322244
rect 378508 322192 378560 322244
rect 518900 322192 518952 322244
rect 346584 321648 346636 321700
rect 346768 321648 346820 321700
rect 259736 321308 259788 321360
rect 259920 321308 259972 321360
rect 249800 320968 249852 321020
rect 314936 320968 314988 321020
rect 350908 320968 350960 321020
rect 401600 320968 401652 321020
rect 178040 320900 178092 320952
rect 297548 320900 297600 320952
rect 378232 320900 378284 320952
rect 523040 320900 523092 320952
rect 131120 320832 131172 320884
rect 286324 320832 286376 320884
rect 287060 320832 287112 320884
rect 287244 320832 287296 320884
rect 389180 320832 389232 320884
rect 565820 320832 565872 320884
rect 3516 320084 3568 320136
rect 233976 320084 234028 320136
rect 252560 319540 252612 319592
rect 305736 319540 305788 319592
rect 350816 319540 350868 319592
rect 405740 319540 405792 319592
rect 200120 319472 200172 319524
rect 303896 319472 303948 319524
rect 357716 319472 357768 319524
rect 432052 319472 432104 319524
rect 84200 319404 84252 319456
rect 276204 319404 276256 319456
rect 381452 319404 381504 319456
rect 532700 319404 532752 319456
rect 197360 318180 197412 318232
rect 302608 318180 302660 318232
rect 355048 318180 355100 318232
rect 419540 318180 419592 318232
rect 184940 318112 184992 318164
rect 299664 318112 299716 318164
rect 361856 318112 361908 318164
rect 448612 318112 448664 318164
rect 93860 318044 93912 318096
rect 279056 318044 279108 318096
rect 303620 318044 303672 318096
rect 327448 318044 327500 318096
rect 382464 318044 382516 318096
rect 539600 318044 539652 318096
rect 218060 316820 218112 316872
rect 307944 316820 307996 316872
rect 349436 316820 349488 316872
rect 398840 316820 398892 316872
rect 193220 316752 193272 316804
rect 301136 316752 301188 316804
rect 356428 316752 356480 316804
rect 423680 316752 423732 316804
rect 60740 316684 60792 316736
rect 263876 316684 263928 316736
rect 264060 316684 264112 316736
rect 338672 316684 338724 316736
rect 349252 316684 349304 316736
rect 385592 316684 385644 316736
rect 550640 316684 550692 316736
rect 270776 316616 270828 316668
rect 211160 315392 211212 315444
rect 306564 315392 306616 315444
rect 360936 315392 360988 315444
rect 430580 315392 430632 315444
rect 128360 315324 128412 315376
rect 287244 315324 287296 315376
rect 365904 315324 365956 315376
rect 466460 315324 466512 315376
rect 66260 315256 66312 315308
rect 272064 315256 272116 315308
rect 386788 315256 386840 315308
rect 554780 315256 554832 315308
rect 229100 314032 229152 314084
rect 310796 314032 310848 314084
rect 195980 313964 196032 314016
rect 302516 313964 302568 314016
rect 368756 313964 368808 314016
rect 481640 313964 481692 314016
rect 57980 313896 58032 313948
rect 270500 313896 270552 313948
rect 343824 313896 343876 313948
rect 372712 313896 372764 313948
rect 386696 313896 386748 313948
rect 557540 313896 557592 313948
rect 282184 313216 282236 313268
rect 580172 313216 580224 313268
rect 223580 312672 223632 312724
rect 309416 312672 309468 312724
rect 135260 312604 135312 312656
rect 287796 312604 287848 312656
rect 44180 312536 44232 312588
rect 266636 312536 266688 312588
rect 353392 312536 353444 312588
rect 416780 312536 416832 312588
rect 236092 311244 236144 311296
rect 312084 311244 312136 311296
rect 347964 311244 348016 311296
rect 389180 311244 389232 311296
rect 202880 311176 202932 311228
rect 303988 311176 304040 311228
rect 357624 311176 357676 311228
rect 434720 311176 434772 311228
rect 4804 311108 4856 311160
rect 256884 311108 256936 311160
rect 388168 311108 388220 311160
rect 561680 311108 561732 311160
rect 209780 309884 209832 309936
rect 305184 309884 305236 309936
rect 350724 309884 350776 309936
rect 402980 309884 403032 309936
rect 147680 309816 147732 309868
rect 291476 309816 291528 309868
rect 364616 309816 364668 309868
rect 459560 309816 459612 309868
rect 77300 309748 77352 309800
rect 273904 309748 273956 309800
rect 388076 309748 388128 309800
rect 564440 309748 564492 309800
rect 227720 308524 227772 308576
rect 309324 308524 309376 308576
rect 143540 308456 143592 308508
rect 289912 308456 289964 308508
rect 352104 308456 352156 308508
rect 409880 308456 409932 308508
rect 18604 308388 18656 308440
rect 258172 308388 258224 308440
rect 389548 308388 389600 308440
rect 567844 308388 567896 308440
rect 245660 307164 245712 307216
rect 313464 307164 313516 307216
rect 179420 307096 179472 307148
rect 298192 307096 298244 307148
rect 356336 307096 356388 307148
rect 427820 307096 427872 307148
rect 75920 307028 75972 307080
rect 274916 307028 274968 307080
rect 345296 307028 345348 307080
rect 378232 307028 378284 307080
rect 390928 307028 390980 307080
rect 575480 307028 575532 307080
rect 2780 306212 2832 306264
rect 4896 306212 4948 306264
rect 247040 305736 247092 305788
rect 314844 305736 314896 305788
rect 353576 305736 353628 305788
rect 415400 305736 415452 305788
rect 139400 305668 139452 305720
rect 288624 305668 288676 305720
rect 367284 305668 367336 305720
rect 473360 305668 473412 305720
rect 40040 305600 40092 305652
rect 264244 305600 264296 305652
rect 339684 305600 339736 305652
rect 353392 305600 353444 305652
rect 378416 305600 378468 305652
rect 521660 305600 521712 305652
rect 201592 304376 201644 304428
rect 303804 304376 303856 304428
rect 143632 304308 143684 304360
rect 289176 304308 289228 304360
rect 354680 304308 354732 304360
rect 423772 304308 423824 304360
rect 88340 304240 88392 304292
rect 277768 304240 277820 304292
rect 372988 304240 373040 304292
rect 495440 304240 495492 304292
rect 219440 303016 219492 303068
rect 307852 303016 307904 303068
rect 146300 302948 146352 303000
rect 291384 302948 291436 303000
rect 357532 302948 357584 303000
rect 433340 302948 433392 303000
rect 27620 302880 27672 302932
rect 262404 302880 262456 302932
rect 377404 302880 377456 302932
rect 509240 302880 509292 302932
rect 230480 301588 230532 301640
rect 310704 301588 310756 301640
rect 150440 301520 150492 301572
rect 291292 301520 291344 301572
rect 359004 301520 359056 301572
rect 437480 301520 437532 301572
rect 22744 301452 22796 301504
rect 259736 301452 259788 301504
rect 378324 301452 378376 301504
rect 520280 301452 520332 301504
rect 153200 300160 153252 300212
rect 292764 300160 292816 300212
rect 358912 300160 358964 300212
rect 440332 300160 440384 300212
rect 110512 300092 110564 300144
rect 283288 300092 283340 300144
rect 381176 300092 381228 300144
rect 531320 300092 531372 300144
rect 567936 299412 567988 299464
rect 579620 299412 579672 299464
rect 157340 298800 157392 298852
rect 292672 298800 292724 298852
rect 360384 298800 360436 298852
rect 444380 298800 444432 298852
rect 26240 298732 26292 298784
rect 261484 298732 261536 298784
rect 385040 298732 385092 298784
rect 552020 298732 552072 298784
rect 255320 297508 255372 297560
rect 316224 297508 316276 297560
rect 126980 297440 127032 297492
rect 285956 297440 286008 297492
rect 361672 297440 361724 297492
rect 451280 297440 451332 297492
rect 102140 297372 102192 297424
rect 280344 297372 280396 297424
rect 390652 297372 390704 297424
rect 572076 297372 572128 297424
rect 165620 296012 165672 296064
rect 295432 296012 295484 296064
rect 363236 296012 363288 296064
rect 455420 296012 455472 296064
rect 35900 295944 35952 295996
rect 265256 295944 265308 295996
rect 365812 295944 365864 295996
rect 470600 295944 470652 295996
rect 176660 294652 176712 294704
rect 297456 294652 297508 294704
rect 363144 294652 363196 294704
rect 458180 294652 458232 294704
rect 20720 294584 20772 294636
rect 261116 294584 261168 294636
rect 296720 294584 296772 294636
rect 325884 294584 325936 294636
rect 371240 294584 371292 294636
rect 490012 294584 490064 294636
rect 3056 293904 3108 293956
rect 221464 293904 221516 293956
rect 369124 293292 369176 293344
rect 465172 293292 465224 293344
rect 215300 293224 215352 293276
rect 306472 293224 306524 293276
rect 375472 293224 375524 293276
rect 506480 293224 506532 293276
rect 299664 292000 299716 292052
rect 327356 292000 327408 292052
rect 183560 291864 183612 291916
rect 299572 291864 299624 291916
rect 367468 291864 367520 291916
rect 476120 291864 476172 291916
rect 29000 291796 29052 291848
rect 263876 291796 263928 291848
rect 342536 291796 342588 291848
rect 367284 291796 367336 291848
rect 379612 291796 379664 291848
rect 524420 291796 524472 291848
rect 190460 290504 190512 290556
rect 301044 290504 301096 290556
rect 370044 290504 370096 290556
rect 484400 290504 484452 290556
rect 114560 290436 114612 290488
rect 283196 290436 283248 290488
rect 383752 290436 383804 290488
rect 542360 290436 542412 290488
rect 193312 289144 193364 289196
rect 302424 289144 302476 289196
rect 16580 289076 16632 289128
rect 256148 289076 256200 289128
rect 369952 289076 370004 289128
rect 488540 289076 488592 289128
rect 129740 287716 129792 287768
rect 287152 287716 287204 287768
rect 60832 287648 60884 287700
rect 269764 287648 269816 287700
rect 345664 287648 345716 287700
rect 371240 287648 371292 287700
rect 371424 287648 371476 287700
rect 491300 287648 491352 287700
rect 208400 286356 208452 286408
rect 305092 286356 305144 286408
rect 96620 286288 96672 286340
rect 278964 286288 279016 286340
rect 372896 286288 372948 286340
rect 498292 286288 498344 286340
rect 307760 285132 307812 285184
rect 328828 285132 328880 285184
rect 222200 284996 222252 285048
rect 308036 284996 308088 285048
rect 78680 284928 78732 284980
rect 274824 284928 274876 284980
rect 343732 284928 343784 284980
rect 374092 284928 374144 284980
rect 374368 284928 374420 284980
rect 502340 284928 502392 284980
rect 226340 283636 226392 283688
rect 309232 283636 309284 283688
rect 89720 283568 89772 283620
rect 277676 283568 277728 283620
rect 374276 283568 374328 283620
rect 506572 283568 506624 283620
rect 133880 282140 133932 282192
rect 287336 282140 287388 282192
rect 376944 282140 376996 282192
rect 516140 282140 516192 282192
rect 233240 280848 233292 280900
rect 310612 280848 310664 280900
rect 64880 280780 64932 280832
rect 268384 280780 268436 280832
rect 381084 280780 381136 280832
rect 534080 280780 534132 280832
rect 240140 279488 240192 279540
rect 311992 279488 312044 279540
rect 8944 279420 8996 279472
rect 256792 279420 256844 279472
rect 346676 279420 346728 279472
rect 382464 279420 382516 279472
rect 382556 279420 382608 279472
rect 538220 279420 538272 279472
rect 314660 278196 314712 278248
rect 330024 278196 330076 278248
rect 251180 278060 251232 278112
rect 315028 278060 315080 278112
rect 7564 277992 7616 278044
rect 256976 277992 257028 278044
rect 346584 277992 346636 278044
rect 385040 277992 385092 278044
rect 385316 277992 385368 278044
rect 547972 277992 548024 278044
rect 151820 276632 151872 276684
rect 291568 276632 291620 276684
rect 386604 276632 386656 276684
rect 556160 276632 556212 276684
rect 162860 275340 162912 275392
rect 294144 275340 294196 275392
rect 81440 275272 81492 275324
rect 276112 275272 276164 275324
rect 387984 275272 388036 275324
rect 563060 275272 563112 275324
rect 167000 273980 167052 274032
rect 295616 273980 295668 274032
rect 99380 273912 99432 273964
rect 280252 273912 280304 273964
rect 389456 273912 389508 273964
rect 569960 273912 570012 273964
rect 431224 273164 431276 273216
rect 579896 273164 579948 273216
rect 169760 272552 169812 272604
rect 296904 272552 296956 272604
rect 106280 272484 106332 272536
rect 281816 272484 281868 272536
rect 353484 272484 353536 272536
rect 414020 272484 414072 272536
rect 173900 271124 173952 271176
rect 296812 271124 296864 271176
rect 347872 271124 347924 271176
rect 390652 271124 390704 271176
rect 390836 271124 390888 271176
rect 574744 271124 574796 271176
rect 180800 269832 180852 269884
rect 298284 269832 298336 269884
rect 354956 269832 355008 269884
rect 420920 269832 420972 269884
rect 63500 269764 63552 269816
rect 271972 269764 272024 269816
rect 341524 269764 341576 269816
rect 354680 269764 354732 269816
rect 385224 269764 385276 269816
rect 549260 269764 549312 269816
rect 185032 268404 185084 268456
rect 298744 268404 298796 268456
rect 70400 268336 70452 268388
rect 273536 268336 273588 268388
rect 360292 268336 360344 268388
rect 445760 268336 445812 268388
rect 3516 267656 3568 267708
rect 232504 267656 232556 267708
rect 234712 266976 234764 267028
rect 310888 266976 310940 267028
rect 361580 266976 361632 267028
rect 452660 266976 452712 267028
rect 187700 265616 187752 265668
rect 300952 265616 301004 265668
rect 363052 265616 363104 265668
rect 456892 265616 456944 265668
rect 191840 264188 191892 264240
rect 301228 264188 301280 264240
rect 364524 264188 364576 264240
rect 463700 264188 463752 264240
rect 198740 262896 198792 262948
rect 302332 262896 302384 262948
rect 41420 262828 41472 262880
rect 266544 262828 266596 262880
rect 367376 262828 367428 262880
rect 473452 262828 473504 262880
rect 135352 261468 135404 261520
rect 288532 261468 288584 261520
rect 368664 261468 368716 261520
rect 477500 261468 477552 261520
rect 241520 260176 241572 260228
rect 313372 260176 313424 260228
rect 52460 260108 52512 260160
rect 269396 260108 269448 260160
rect 369860 260108 369912 260160
rect 485780 260108 485832 260160
rect 407856 259360 407908 259412
rect 579804 259360 579856 259412
rect 138020 258680 138072 258732
rect 288716 258680 288768 258732
rect 354864 258680 354916 258732
rect 418160 258680 418212 258732
rect 144920 257320 144972 257372
rect 290096 257320 290148 257372
rect 371332 257320 371384 257372
rect 492680 257320 492732 257372
rect 151912 255960 151964 256012
rect 292948 255960 293000 256012
rect 372804 255960 372856 256012
rect 499580 255960 499632 256012
rect 3148 255212 3200 255264
rect 14556 255212 14608 255264
rect 69020 254532 69072 254584
rect 271236 254532 271288 254584
rect 374184 254532 374236 254584
rect 503720 254532 503772 254584
rect 82820 253172 82872 253224
rect 275284 253172 275336 253224
rect 375380 253172 375432 253224
rect 510620 253172 510672 253224
rect 100760 251812 100812 251864
rect 279424 251812 279476 251864
rect 376852 251812 376904 251864
rect 517520 251812 517572 251864
rect 118700 250452 118752 250504
rect 284576 250452 284628 250504
rect 379520 250452 379572 250504
rect 528560 250452 528612 250504
rect 2780 249024 2832 249076
rect 256056 249024 256108 249076
rect 380992 249024 381044 249076
rect 535460 249024 535512 249076
rect 48320 247664 48372 247716
rect 267924 247664 267976 247716
rect 383660 247664 383712 247716
rect 546500 247664 546552 247716
rect 59360 246304 59412 246356
rect 270592 246304 270644 246356
rect 385132 246304 385184 246356
rect 553400 246304 553452 246356
rect 422944 245556 422996 245608
rect 580172 245556 580224 245608
rect 62120 244876 62172 244928
rect 270868 244876 270920 244928
rect 354772 244876 354824 244928
rect 422300 244876 422352 244928
rect 73160 243516 73212 243568
rect 273444 243516 273496 243568
rect 387892 243516 387944 243568
rect 560300 243516 560352 243568
rect 80060 242156 80112 242208
rect 274732 242156 274784 242208
rect 389364 242156 389416 242208
rect 567200 242156 567252 242208
rect 3516 241408 3568 241460
rect 220084 241408 220136 241460
rect 237472 240728 237524 240780
rect 312176 240728 312228 240780
rect 393964 240728 394016 240780
rect 578240 240728 578292 240780
rect 93952 239368 94004 239420
rect 278872 239368 278924 239420
rect 111800 238008 111852 238060
rect 283104 238008 283156 238060
rect 115940 236648 115992 236700
rect 283012 236648 283064 236700
rect 30380 235220 30432 235272
rect 263784 235220 263836 235272
rect 39304 233860 39356 233912
rect 265164 233860 265216 233912
rect 395436 233180 395488 233232
rect 580172 233180 580224 233232
rect 44272 232500 44324 232552
rect 266452 232500 266504 232552
rect 49700 231072 49752 231124
rect 267832 231072 267884 231124
rect 52552 229712 52604 229764
rect 269304 229712 269356 229764
rect 56600 228352 56652 228404
rect 269212 228352 269264 228404
rect 67640 226992 67692 227044
rect 272156 226992 272208 227044
rect 74540 225564 74592 225616
rect 273352 225564 273404 225616
rect 13820 224204 13872 224256
rect 259644 224204 259696 224256
rect 158720 222844 158772 222896
rect 293316 222844 293368 222896
rect 85672 221416 85724 221468
rect 276296 221416 276348 221468
rect 92480 220056 92532 220108
rect 277584 220056 277636 220108
rect 432604 219376 432656 219428
rect 579896 219376 579948 219428
rect 102232 218696 102284 218748
rect 280436 218696 280488 218748
rect 3332 215228 3384 215280
rect 18696 215228 18748 215280
rect 17960 214548 18012 214600
rect 261024 214548 261076 214600
rect 421564 206932 421616 206984
rect 580172 206932 580224 206984
rect 3056 202784 3108 202836
rect 90364 202784 90416 202836
rect 428464 193128 428516 193180
rect 580172 193128 580224 193180
rect 3516 188980 3568 189032
rect 217324 188980 217376 189032
rect 216680 188300 216732 188352
rect 306656 188300 306708 188352
rect 386512 182792 386564 182844
rect 558920 182792 558972 182844
rect 405004 179324 405056 179376
rect 579988 179324 580040 179376
rect 350632 178644 350684 178696
rect 404360 178644 404412 178696
rect 390744 171776 390796 171828
rect 574100 171776 574152 171828
rect 418804 166948 418856 167000
rect 580172 166948 580224 167000
rect 251272 166268 251324 166320
rect 314752 166268 314804 166320
rect 3240 164160 3292 164212
rect 229744 164160 229796 164212
rect 554044 153144 554096 153196
rect 579804 153144 579856 153196
rect 346492 140020 346544 140072
rect 386512 140020 386564 140072
rect 3516 137232 3568 137284
rect 414112 137232 414164 137284
rect 417424 126896 417476 126948
rect 580172 126896 580224 126948
rect 427084 113092 427136 113144
rect 580172 113092 580224 113144
rect 3148 111732 3200 111784
rect 228364 111732 228416 111784
rect 250444 100648 250496 100700
rect 580172 100648 580224 100700
rect 389272 90312 389324 90364
rect 570604 90312 570656 90364
rect 414664 86912 414716 86964
rect 580172 86912 580224 86964
rect 350540 86232 350592 86284
rect 400220 86232 400272 86284
rect 3424 85484 3476 85536
rect 400864 85484 400916 85536
rect 424324 73108 424376 73160
rect 579988 73108 580040 73160
rect 3424 71680 3476 71732
rect 225604 71680 225656 71732
rect 246304 60664 246356 60716
rect 580172 60664 580224 60716
rect 127072 51688 127124 51740
rect 285864 51688 285916 51740
rect 285956 51688 286008 51740
rect 323124 51688 323176 51740
rect 113180 48968 113232 49020
rect 282920 48968 282972 49020
rect 345204 47676 345256 47728
rect 382556 47676 382608 47728
rect 95240 47540 95292 47592
rect 279148 47540 279200 47592
rect 382372 47540 382424 47592
rect 540980 47540 541032 47592
rect 238024 46180 238076 46232
rect 580356 46180 580408 46232
rect 122840 43392 122892 43444
rect 285772 43392 285824 43444
rect 77392 42032 77444 42084
rect 275008 42032 275060 42084
rect 9680 40672 9732 40724
rect 257436 40672 257488 40724
rect 69112 39312 69164 39364
rect 271144 39312 271196 39364
rect 140780 37884 140832 37936
rect 289084 37884 289136 37936
rect 55220 36524 55272 36576
rect 269488 36524 269540 36576
rect 160192 35164 160244 35216
rect 293224 35164 293276 35216
rect 244280 33736 244332 33788
rect 313648 33736 313700 33788
rect 3424 33056 3476 33108
rect 224224 33056 224276 33108
rect 237380 33056 237432 33108
rect 580172 33056 580224 33108
rect 226432 31016 226484 31068
rect 309508 31016 309560 31068
rect 212540 29588 212592 29640
rect 302884 29588 302936 29640
rect 352012 29588 352064 29640
rect 407212 29588 407264 29640
rect 209872 28228 209924 28280
rect 305276 28228 305328 28280
rect 349344 28228 349396 28280
rect 397460 28228 397512 28280
rect 194600 26868 194652 26920
rect 302240 26868 302292 26920
rect 347780 26868 347832 26920
rect 393320 26868 393372 26920
rect 186320 25508 186372 25560
rect 299848 25508 299900 25560
rect 343640 25508 343692 25560
rect 375380 25508 375432 25560
rect 176752 24080 176804 24132
rect 296168 24080 296220 24132
rect 341064 24080 341116 24132
rect 361580 24080 361632 24132
rect 382280 24080 382332 24132
rect 539692 24080 539744 24132
rect 154580 22720 154632 22772
rect 291844 22720 291896 22772
rect 292580 22720 292632 22772
rect 324504 22720 324556 22772
rect 342444 22720 342496 22772
rect 368664 22720 368716 22772
rect 380900 22720 380952 22772
rect 531412 22720 531464 22772
rect 204260 21360 204312 21412
rect 303712 21360 303764 21412
rect 310520 21360 310572 21412
rect 328736 21360 328788 21412
rect 337108 21360 337160 21412
rect 346492 21360 346544 21412
rect 376760 21360 376812 21412
rect 514760 21360 514812 21412
rect 3424 20612 3476 20664
rect 413376 20612 413428 20664
rect 269120 18640 269172 18692
rect 319076 18640 319128 18692
rect 172520 18572 172572 18624
rect 296076 18572 296128 18624
rect 299480 18572 299532 18624
rect 323676 18572 323728 18624
rect 368572 18572 368624 18624
rect 481732 18572 481784 18624
rect 259644 17280 259696 17332
rect 317604 17280 317656 17332
rect 349160 17280 349212 17332
rect 398932 17280 398984 17332
rect 118792 17212 118844 17264
rect 284484 17212 284536 17264
rect 295340 17212 295392 17264
rect 324964 17212 325016 17264
rect 387800 17212 387852 17264
rect 564532 17212 564584 17264
rect 109040 16056 109092 16108
rect 281632 16056 281684 16108
rect 105728 15988 105780 16040
rect 281724 15988 281776 16040
rect 91560 15920 91612 15972
rect 277400 15920 277452 15972
rect 282000 15920 282052 15972
rect 304264 15920 304316 15972
rect 345112 15920 345164 15972
rect 379520 15920 379572 15972
rect 87512 15852 87564 15904
rect 277492 15852 277544 15904
rect 279056 15852 279108 15904
rect 316684 15852 316736 15904
rect 372620 15852 372672 15904
rect 497096 15852 497148 15904
rect 273352 14560 273404 14612
rect 320364 14560 320416 14612
rect 122288 14492 122340 14544
rect 284392 14492 284444 14544
rect 108120 14424 108172 14476
rect 281908 14424 281960 14476
rect 284576 14424 284628 14476
rect 305644 14424 305696 14476
rect 306380 14424 306432 14476
rect 328644 14424 328696 14476
rect 339592 14424 339644 14476
rect 357532 14424 357584 14476
rect 378140 14424 378192 14476
rect 523776 14424 523828 14476
rect 278320 13200 278372 13252
rect 300124 13200 300176 13252
rect 283104 13132 283156 13184
rect 307024 13132 307076 13184
rect 346400 13132 346452 13184
rect 387800 13132 387852 13184
rect 137192 13064 137244 13116
rect 287704 13064 287756 13116
rect 303160 13064 303212 13116
rect 327264 13064 327316 13116
rect 386420 13064 386472 13116
rect 556896 13064 556948 13116
rect 143540 11772 143592 11824
rect 144736 11772 144788 11824
rect 160100 11772 160152 11824
rect 161296 11772 161348 11824
rect 184940 11772 184992 11824
rect 186136 11772 186188 11824
rect 234620 11772 234672 11824
rect 235816 11772 235868 11824
rect 242900 11772 242952 11824
rect 244096 11772 244148 11824
rect 274824 11772 274876 11824
rect 320272 11772 320324 11824
rect 351920 11772 351972 11824
rect 411904 11772 411956 11824
rect 51080 11704 51132 11756
rect 257344 11704 257396 11756
rect 265164 11704 265216 11756
rect 318984 11704 319036 11756
rect 340972 11704 341024 11756
rect 363512 11704 363564 11756
rect 407764 11704 407816 11756
rect 537208 11704 537260 11756
rect 309876 10480 309928 10532
rect 328552 10480 328604 10532
rect 270776 10412 270828 10464
rect 309784 10412 309836 10464
rect 280712 10344 280764 10396
rect 321652 10344 321704 10396
rect 72608 10276 72660 10328
rect 273628 10276 273680 10328
rect 276020 10276 276072 10328
rect 320456 10276 320508 10328
rect 342352 10276 342404 10328
rect 370136 10276 370188 10328
rect 399484 10276 399536 10328
rect 515496 10276 515548 10328
rect 209688 9596 209740 9648
rect 210976 9596 211028 9648
rect 359464 9596 359516 9648
rect 361120 9596 361172 9648
rect 261760 9052 261812 9104
rect 311164 9052 311216 9104
rect 266544 8984 266596 9036
rect 318892 8984 318944 9036
rect 132960 8916 133012 8968
rect 243544 8916 243596 8968
rect 264152 8916 264204 8968
rect 317512 8916 317564 8968
rect 320916 8916 320968 8968
rect 331496 8916 331548 8968
rect 340880 8916 340932 8968
rect 359924 8916 359976 8968
rect 370504 8916 370556 8968
rect 393044 8916 393096 8968
rect 410524 8916 410576 8968
rect 501788 8916 501840 8968
rect 360844 8372 360896 8424
rect 365812 8372 365864 8424
rect 292580 7760 292632 7812
rect 324412 7760 324464 7812
rect 260656 7692 260708 7744
rect 301504 7692 301556 7744
rect 218152 7624 218204 7676
rect 247684 7624 247736 7676
rect 277124 7624 277176 7676
rect 321744 7624 321796 7676
rect 338396 7624 338448 7676
rect 349160 7624 349212 7676
rect 33600 7556 33652 7608
rect 233884 7556 233936 7608
rect 268844 7556 268896 7608
rect 319168 7556 319220 7608
rect 324412 7556 324464 7608
rect 332968 7556 333020 7608
rect 345020 7556 345072 7608
rect 381176 7556 381228 7608
rect 395344 7556 395396 7608
rect 487620 7556 487672 7608
rect 236000 6808 236052 6860
rect 580172 6808 580224 6860
rect 288992 6264 289044 6316
rect 297364 6264 297416 6316
rect 262956 6196 263008 6248
rect 317696 6196 317748 6248
rect 169576 6128 169628 6180
rect 242164 6128 242216 6180
rect 258264 6128 258316 6180
rect 315304 6128 315356 6180
rect 318524 6128 318576 6180
rect 327724 6128 327776 6180
rect 339500 6128 339552 6180
rect 358728 6128 358780 6180
rect 267740 4972 267792 5024
rect 295984 4972 296036 5024
rect 313832 4972 313884 5024
rect 320824 4972 320876 5024
rect 290188 4904 290240 4956
rect 323584 4904 323636 4956
rect 336924 4904 336976 4956
rect 345756 4904 345808 4956
rect 272432 4836 272484 4888
rect 318064 4836 318116 4888
rect 338304 4836 338356 4888
rect 352840 4836 352892 4888
rect 353300 4836 353352 4888
rect 415492 4836 415544 4888
rect 168380 4768 168432 4820
rect 255964 4768 256016 4820
rect 257068 4768 257120 4820
rect 313924 4768 313976 4820
rect 342260 4768 342312 4820
rect 363604 4768 363656 4820
rect 364616 4768 364668 4820
rect 371884 4768 371936 4820
rect 377680 4768 377732 4820
rect 396724 4768 396776 4820
rect 484032 4768 484084 4820
rect 367008 4700 367060 4752
rect 378784 4496 378836 4548
rect 384764 4496 384816 4548
rect 135260 4156 135312 4208
rect 136456 4156 136508 4208
rect 218060 4156 218112 4208
rect 219256 4156 219308 4208
rect 43076 4088 43128 4140
rect 258448 4156 258500 4208
rect 317328 4156 317380 4208
rect 322204 4156 322256 4208
rect 337016 4156 337068 4208
rect 342168 4156 342220 4208
rect 319720 4088 319772 4140
rect 331404 4088 331456 4140
rect 358820 4088 358872 4140
rect 440240 4088 440292 4140
rect 2872 4020 2924 4072
rect 8944 4020 8996 4072
rect 39580 4020 39632 4072
rect 265072 4020 265124 4072
rect 316224 4020 316276 4072
rect 330116 4020 330168 4072
rect 360200 4020 360252 4072
rect 447416 4020 447468 4072
rect 35992 3952 36044 4004
rect 264980 3952 265032 4004
rect 312636 3952 312688 4004
rect 329932 3952 329984 4004
rect 362960 3952 363012 4004
rect 454500 3952 454552 4004
rect 32404 3884 32456 3936
rect 263968 3884 264020 3936
rect 309048 3884 309100 3936
rect 328460 3884 328512 3936
rect 364340 3884 364392 3936
rect 461584 3884 461636 3936
rect 28908 3816 28960 3868
rect 263692 3816 263744 3868
rect 305552 3816 305604 3868
rect 327172 3816 327224 3868
rect 364432 3816 364484 3868
rect 465172 3816 465224 3868
rect 574744 3816 574796 3868
rect 577412 3816 577464 3868
rect 25320 3748 25372 3800
rect 262312 3748 262364 3800
rect 301964 3748 302016 3800
rect 327080 3748 327132 3800
rect 328000 3748 328052 3800
rect 332692 3748 332744 3800
rect 335452 3748 335504 3800
rect 340972 3748 341024 3800
rect 365720 3748 365772 3800
rect 468668 3748 468720 3800
rect 6460 3680 6512 3732
rect 10324 3680 10376 3732
rect 13544 3680 13596 3732
rect 22744 3680 22796 3732
rect 24216 3680 24268 3732
rect 258080 3680 258132 3732
rect 20628 3612 20680 3664
rect 261208 3680 261260 3732
rect 298468 3680 298520 3732
rect 325976 3680 326028 3732
rect 331588 3680 331640 3732
rect 334072 3680 334124 3732
rect 335728 3680 335780 3732
rect 339868 3680 339920 3732
rect 367100 3680 367152 3732
rect 472256 3680 472308 3732
rect 8760 3544 8812 3596
rect 18604 3544 18656 3596
rect 19432 3544 19484 3596
rect 260932 3612 260984 3664
rect 294880 3612 294932 3664
rect 325792 3612 325844 3664
rect 332692 3612 332744 3664
rect 334164 3612 334216 3664
rect 335636 3612 335688 3664
rect 338672 3612 338724 3664
rect 367192 3612 367244 3664
rect 475752 3612 475804 3664
rect 258448 3544 258500 3596
rect 266728 3544 266780 3596
rect 285680 3544 285732 3596
rect 286048 3544 286100 3596
rect 291384 3544 291436 3596
rect 7656 3476 7708 3528
rect 13084 3476 13136 3528
rect 15936 3476 15988 3528
rect 259368 3476 259420 3528
rect 323308 3544 323360 3596
rect 331312 3544 331364 3596
rect 333980 3544 334032 3596
rect 334716 3544 334768 3596
rect 335544 3544 335596 3596
rect 337476 3544 337528 3596
rect 356152 3544 356204 3596
rect 324596 3476 324648 3528
rect 326804 3476 326856 3528
rect 332876 3476 332928 3528
rect 338120 3476 338172 3528
rect 348056 3476 348108 3528
rect 349252 3476 349304 3528
rect 350448 3476 350500 3528
rect 1676 3408 1728 3460
rect 7564 3408 7616 3460
rect 11152 3408 11204 3460
rect 259828 3408 259880 3460
rect 284300 3408 284352 3460
rect 323032 3408 323084 3460
rect 325608 3408 325660 3460
rect 332600 3408 332652 3460
rect 338212 3408 338264 3460
rect 351644 3408 351696 3460
rect 38384 3340 38436 3392
rect 39304 3340 39356 3392
rect 46664 3340 46716 3392
rect 268108 3340 268160 3392
rect 322112 3340 322164 3392
rect 331496 3340 331548 3392
rect 60740 3272 60792 3324
rect 61660 3272 61712 3324
rect 85580 3272 85632 3324
rect 86500 3272 86552 3324
rect 121092 3272 121144 3324
rect 284668 3272 284720 3324
rect 287796 3272 287848 3324
rect 323216 3272 323268 3324
rect 382464 3544 382516 3596
rect 383568 3544 383620 3596
rect 392124 3544 392176 3596
rect 581000 3544 581052 3596
rect 368480 3476 368532 3528
rect 479340 3476 479392 3528
rect 489920 3476 489972 3528
rect 490748 3476 490800 3528
rect 506480 3476 506532 3528
rect 507308 3476 507360 3528
rect 539600 3476 539652 3528
rect 540428 3476 540480 3528
rect 564440 3476 564492 3528
rect 565268 3476 565320 3528
rect 567844 3476 567896 3528
rect 569132 3476 569184 3528
rect 570604 3476 570656 3528
rect 571524 3476 571576 3528
rect 571984 3476 572036 3528
rect 572720 3476 572772 3528
rect 374092 3408 374144 3460
rect 375288 3408 375340 3460
rect 390560 3408 390612 3460
rect 391848 3408 391900 3460
rect 391940 3408 391992 3460
rect 582196 3408 582248 3460
rect 357440 3340 357492 3392
rect 433248 3340 433300 3392
rect 440332 3340 440384 3392
rect 441528 3340 441580 3392
rect 448612 3340 448664 3392
rect 449808 3340 449860 3392
rect 572076 3340 572128 3392
rect 573916 3340 573968 3392
rect 124680 3204 124732 3256
rect 285680 3204 285732 3256
rect 329196 3204 329248 3256
rect 332784 3204 332836 3256
rect 356428 3204 356480 3256
rect 258080 3136 258132 3188
rect 262588 3136 262640 3188
rect 330392 3136 330444 3188
rect 334348 3136 334400 3188
rect 398932 3136 398984 3188
rect 400128 3136 400180 3188
rect 407212 3136 407264 3188
rect 408408 3136 408460 3188
rect 572 3068 624 3120
rect 4804 3068 4856 3120
rect 23020 3068 23072 3120
rect 25504 3068 25556 3120
rect 415400 3204 415452 3256
rect 416688 3204 416740 3256
rect 423680 3272 423732 3324
rect 424968 3272 425020 3324
rect 429660 3136 429712 3188
rect 426164 3068 426216 3120
rect 12348 3000 12400 3052
rect 14464 3000 14516 3052
rect 336832 3000 336884 3052
rect 344560 3000 344612 3052
rect 336740 2932 336792 2984
rect 343364 2932 343416 2984
rect 456800 1640 456852 1692
rect 458088 1640 458140 1692
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 700330 8156 703520
rect 24320 700398 24348 703520
rect 24308 700392 24360 700398
rect 24308 700334 24360 700340
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3330 619168 3386 619177
rect 3330 619103 3386 619112
rect 3344 618322 3372 619103
rect 3332 618316 3384 618322
rect 3332 618258 3384 618264
rect 3330 606112 3386 606121
rect 3330 606047 3386 606056
rect 3344 605878 3372 606047
rect 3332 605872 3384 605878
rect 3332 605814 3384 605820
rect 3054 566944 3110 566953
rect 3054 566879 3110 566888
rect 3068 565894 3096 566879
rect 3056 565888 3108 565894
rect 3056 565830 3108 565836
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 3330 514856 3386 514865
rect 3330 514791 3332 514800
rect 3384 514791 3386 514800
rect 3332 514762 3384 514768
rect 3238 501800 3294 501809
rect 3238 501735 3294 501744
rect 3252 501022 3280 501735
rect 3240 501016 3292 501022
rect 3240 500958 3292 500964
rect 3436 460193 3464 684247
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3514 658200 3570 658209
rect 3514 658135 3570 658144
rect 3528 656946 3556 658135
rect 3516 656940 3568 656946
rect 3516 656882 3568 656888
rect 3514 632088 3570 632097
rect 3514 632023 3570 632032
rect 3528 465746 3556 632023
rect 3606 580000 3662 580009
rect 3606 579935 3662 579944
rect 3620 465882 3648 579935
rect 3698 527912 3754 527921
rect 3698 527847 3754 527856
rect 3712 466018 3740 527847
rect 3882 475688 3938 475697
rect 3882 475623 3938 475632
rect 3712 465990 3832 466018
rect 3620 465854 3740 465882
rect 3528 465718 3648 465746
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3528 462398 3556 462567
rect 3516 462392 3568 462398
rect 3516 462334 3568 462340
rect 3620 460426 3648 465718
rect 3608 460420 3660 460426
rect 3608 460362 3660 460368
rect 3712 460358 3740 465854
rect 3700 460352 3752 460358
rect 3700 460294 3752 460300
rect 3804 460290 3832 465990
rect 3792 460284 3844 460290
rect 3792 460226 3844 460232
rect 3896 460222 3924 475623
rect 40052 474026 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 40040 474020 40092 474026
rect 40040 473962 40092 473968
rect 13084 463752 13136 463758
rect 13084 463694 13136 463700
rect 3884 460216 3936 460222
rect 3422 460184 3478 460193
rect 3884 460158 3936 460164
rect 3422 460119 3478 460128
rect 3424 458244 3476 458250
rect 3424 458186 3476 458192
rect 3436 423609 3464 458186
rect 3516 457496 3568 457502
rect 3516 457438 3568 457444
rect 3528 449585 3556 457438
rect 3514 449576 3570 449585
rect 3514 449511 3570 449520
rect 3422 423600 3478 423609
rect 3422 423535 3478 423544
rect 3424 411256 3476 411262
rect 3424 411198 3476 411204
rect 3436 410553 3464 411198
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 3240 398812 3292 398818
rect 3240 398754 3292 398760
rect 3252 397497 3280 398754
rect 3238 397488 3294 397497
rect 3238 397423 3294 397432
rect 3240 372564 3292 372570
rect 3240 372506 3292 372512
rect 3252 371385 3280 372506
rect 3238 371376 3294 371385
rect 3238 371311 3294 371320
rect 3332 358760 3384 358766
rect 3332 358702 3384 358708
rect 3344 358465 3372 358702
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 13096 346390 13124 463694
rect 18696 460964 18748 460970
rect 18696 460906 18748 460912
rect 3148 346384 3200 346390
rect 3148 346326 3200 346332
rect 13084 346384 13136 346390
rect 13084 346326 13136 346332
rect 3160 345409 3188 346326
rect 3146 345400 3202 345409
rect 3146 345335 3202 345344
rect 3422 337376 3478 337385
rect 3422 337311 3478 337320
rect 2780 306264 2832 306270
rect 2778 306232 2780 306241
rect 2832 306232 2834 306241
rect 2778 306167 2834 306176
rect 3056 293956 3108 293962
rect 3056 293898 3108 293904
rect 3068 293185 3096 293898
rect 3054 293176 3110 293185
rect 3054 293111 3110 293120
rect 3148 255264 3200 255270
rect 3148 255206 3200 255212
rect 3160 254153 3188 255206
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 2780 249076 2832 249082
rect 2780 249018 2832 249024
rect 2792 16574 2820 249018
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3056 202836 3108 202842
rect 3056 202778 3108 202784
rect 3068 201929 3096 202778
rect 3054 201920 3110 201929
rect 3054 201855 3110 201864
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3436 136785 3464 337311
rect 10324 336048 10376 336054
rect 10324 335990 10376 335996
rect 4894 331800 4950 331809
rect 4894 331735 4950 331744
rect 3516 320136 3568 320142
rect 3516 320078 3568 320084
rect 3528 319297 3556 320078
rect 3514 319288 3570 319297
rect 3514 319223 3570 319232
rect 4804 311160 4856 311166
rect 4804 311102 4856 311108
rect 3516 267708 3568 267714
rect 3516 267650 3568 267656
rect 3528 267209 3556 267650
rect 3514 267200 3570 267209
rect 3514 267135 3570 267144
rect 3516 241460 3568 241466
rect 3516 241402 3568 241408
rect 3528 241097 3556 241402
rect 3514 241088 3570 241097
rect 3514 241023 3570 241032
rect 3516 189032 3568 189038
rect 3516 188974 3568 188980
rect 3528 188873 3556 188974
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 3516 137284 3568 137290
rect 3516 137226 3568 137232
rect 3422 136776 3478 136785
rect 3422 136711 3478 136720
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 3424 85536 3476 85542
rect 3424 85478 3476 85484
rect 3436 84697 3464 85478
rect 3422 84688 3478 84697
rect 3422 84623 3478 84632
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3424 33108 3476 33114
rect 3424 33050 3476 33056
rect 3436 32473 3464 33050
rect 3422 32464 3478 32473
rect 3422 32399 3478 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 2792 16546 3464 16574
rect 2872 4072 2924 4078
rect 2872 4014 2924 4020
rect 1676 3460 1728 3466
rect 1676 3402 1728 3408
rect 572 3120 624 3126
rect 572 3062 624 3068
rect 584 480 612 3062
rect 1688 480 1716 3402
rect 2884 480 2912 4014
rect 3436 490 3464 16546
rect 3528 6497 3556 137226
rect 3514 6488 3570 6497
rect 3514 6423 3570 6432
rect 4816 3126 4844 311102
rect 4908 306270 4936 331735
rect 4896 306264 4948 306270
rect 4896 306206 4948 306212
rect 8944 279472 8996 279478
rect 8944 279414 8996 279420
rect 7564 278044 7616 278050
rect 7564 277986 7616 277992
rect 6460 3732 6512 3738
rect 6460 3674 6512 3680
rect 5262 3360 5318 3369
rect 5262 3295 5318 3304
rect 4804 3120 4856 3126
rect 4804 3062 4856 3068
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3436 462 3648 490
rect 5276 480 5304 3295
rect 6472 480 6500 3674
rect 7576 3466 7604 277986
rect 8956 4078 8984 279414
rect 9680 40724 9732 40730
rect 9680 40666 9732 40672
rect 8944 4072 8996 4078
rect 8944 4014 8996 4020
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7564 3460 7616 3466
rect 7564 3402 7616 3408
rect 7668 480 7696 3470
rect 8772 480 8800 3538
rect 3620 354 3648 462
rect 4038 354 4150 480
rect 3620 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 40666
rect 10336 3738 10364 335990
rect 14464 334620 14516 334626
rect 14464 334562 14516 334568
rect 13084 333260 13136 333266
rect 13084 333202 13136 333208
rect 10324 3732 10376 3738
rect 10324 3674 10376 3680
rect 13096 3534 13124 333202
rect 13820 224256 13872 224262
rect 13820 224198 13872 224204
rect 13832 16574 13860 224198
rect 13832 16546 14320 16574
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11164 480 11192 3402
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 12360 480 12388 2994
rect 13556 480 13584 3674
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 14476 3058 14504 334562
rect 14554 330440 14610 330449
rect 14554 330375 14610 330384
rect 14568 255270 14596 330375
rect 18604 308440 18656 308446
rect 18604 308382 18656 308388
rect 16580 289128 16632 289134
rect 16580 289070 16632 289076
rect 14556 255264 14608 255270
rect 14556 255206 14608 255212
rect 16592 16574 16620 289070
rect 17960 214600 18012 214606
rect 17960 214542 18012 214548
rect 16592 16546 17080 16574
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 14464 3052 14516 3058
rect 14464 2994 14516 3000
rect 15948 480 15976 3470
rect 17052 480 17080 16546
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 214542
rect 18616 3602 18644 308382
rect 18708 215286 18736 460906
rect 71792 460494 71820 702986
rect 89180 700466 89208 703520
rect 89168 700460 89220 700466
rect 89168 700402 89220 700408
rect 105464 699718 105492 703520
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106924 699712 106976 699718
rect 106924 699654 106976 699660
rect 106936 469878 106964 699654
rect 106924 469872 106976 469878
rect 106924 469814 106976 469820
rect 136652 460698 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 700534 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 169772 702406 170352 702434
rect 154120 700528 154172 700534
rect 154120 700470 154172 700476
rect 169772 468518 169800 702406
rect 169760 468512 169812 468518
rect 169760 468454 169812 468460
rect 201512 460902 201540 702986
rect 218992 700602 219020 703520
rect 218980 700596 219032 700602
rect 218980 700538 219032 700544
rect 234632 467158 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 697610 267688 703520
rect 283852 700738 283880 703520
rect 283840 700732 283892 700738
rect 283840 700674 283892 700680
rect 300136 700058 300164 703520
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 322940 700800 322992 700806
rect 322940 700742 322992 700748
rect 318800 700664 318852 700670
rect 318800 700606 318852 700612
rect 300124 700052 300176 700058
rect 300124 699994 300176 700000
rect 301504 700052 301556 700058
rect 301504 699994 301556 700000
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 234620 467152 234672 467158
rect 234620 467094 234672 467100
rect 215944 464024 215996 464030
rect 215944 463966 215996 463972
rect 201500 460896 201552 460902
rect 201500 460838 201552 460844
rect 136640 460692 136692 460698
rect 136640 460634 136692 460640
rect 71780 460488 71832 460494
rect 71780 460430 71832 460436
rect 215956 358766 215984 463966
rect 220084 463956 220136 463962
rect 220084 463898 220136 463904
rect 217324 463888 217376 463894
rect 217324 463830 217376 463836
rect 215944 358760 215996 358766
rect 215944 358702 215996 358708
rect 117320 336184 117372 336190
rect 117320 336126 117372 336132
rect 110420 336116 110472 336122
rect 110420 336058 110472 336064
rect 98000 331900 98052 331906
rect 98000 331842 98052 331848
rect 90362 329080 90418 329089
rect 90362 329015 90418 329024
rect 85580 327752 85632 327758
rect 85580 327694 85632 327700
rect 53840 326392 53892 326398
rect 53840 326334 53892 326340
rect 46940 324964 46992 324970
rect 46940 324906 46992 324912
rect 25504 323604 25556 323610
rect 25504 323546 25556 323552
rect 22744 301504 22796 301510
rect 22744 301446 22796 301452
rect 20720 294636 20772 294642
rect 20720 294578 20772 294584
rect 18696 215280 18748 215286
rect 18696 215222 18748 215228
rect 20732 16574 20760 294578
rect 20732 16546 21864 16574
rect 20628 3664 20680 3670
rect 20628 3606 20680 3612
rect 18604 3596 18656 3602
rect 18604 3538 18656 3544
rect 19432 3596 19484 3602
rect 19432 3538 19484 3544
rect 19444 480 19472 3538
rect 20640 480 20668 3606
rect 21836 480 21864 16546
rect 22756 3738 22784 301446
rect 25320 3800 25372 3806
rect 25320 3742 25372 3748
rect 22744 3732 22796 3738
rect 22744 3674 22796 3680
rect 24216 3732 24268 3738
rect 24216 3674 24268 3680
rect 23020 3120 23072 3126
rect 23020 3062 23072 3068
rect 23032 480 23060 3062
rect 24228 480 24256 3674
rect 25332 480 25360 3742
rect 25516 3126 25544 323546
rect 34520 322244 34572 322250
rect 34520 322186 34572 322192
rect 27620 302932 27672 302938
rect 27620 302874 27672 302880
rect 26240 298784 26292 298790
rect 26240 298726 26292 298732
rect 25504 3120 25556 3126
rect 25504 3062 25556 3068
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 298726
rect 27632 16574 27660 302874
rect 29000 291848 29052 291854
rect 29000 291790 29052 291796
rect 29012 16574 29040 291790
rect 30380 235272 30432 235278
rect 30380 235214 30432 235220
rect 30392 16574 30420 235214
rect 27632 16546 27752 16574
rect 29012 16546 30144 16574
rect 30392 16546 30880 16574
rect 27724 480 27752 16546
rect 28908 3868 28960 3874
rect 28908 3810 28960 3816
rect 28920 480 28948 3810
rect 30116 480 30144 16546
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 33600 7608 33652 7614
rect 33600 7550 33652 7556
rect 32404 3936 32456 3942
rect 32404 3878 32456 3884
rect 32416 480 32444 3878
rect 33612 480 33640 7550
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31270 -960 31382 326
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34532 354 34560 322186
rect 44180 312588 44232 312594
rect 44180 312530 44232 312536
rect 40040 305652 40092 305658
rect 40040 305594 40092 305600
rect 35900 295996 35952 296002
rect 35900 295938 35952 295944
rect 35912 16574 35940 295938
rect 39304 233912 39356 233918
rect 39304 233854 39356 233860
rect 35912 16546 36768 16574
rect 35992 4004 36044 4010
rect 35992 3946 36044 3952
rect 36004 480 36032 3946
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 39316 3398 39344 233854
rect 40052 16574 40080 305594
rect 41420 262880 41472 262886
rect 41420 262822 41472 262828
rect 41432 16574 41460 262822
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 39580 4072 39632 4078
rect 39580 4014 39632 4020
rect 38384 3392 38436 3398
rect 38384 3334 38436 3340
rect 39304 3392 39356 3398
rect 39304 3334 39356 3340
rect 38396 480 38424 3334
rect 39592 480 39620 4014
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40236 354 40264 16546
rect 41892 480 41920 16546
rect 44192 6914 44220 312530
rect 44272 232552 44324 232558
rect 44272 232494 44324 232500
rect 44284 16574 44312 232494
rect 46952 16574 46980 324906
rect 52460 260160 52512 260166
rect 52460 260102 52512 260108
rect 48320 247716 48372 247722
rect 48320 247658 48372 247664
rect 48332 16574 48360 247658
rect 49700 231124 49752 231130
rect 49700 231066 49752 231072
rect 49712 16574 49740 231066
rect 44284 16546 45048 16574
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 44192 6886 44312 6914
rect 43076 4140 43128 4146
rect 43076 4082 43128 4088
rect 43088 480 43116 4082
rect 44284 480 44312 6886
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 46664 3392 46716 3398
rect 46664 3334 46716 3340
rect 46676 480 46704 3334
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 51080 11756 51132 11762
rect 51080 11698 51132 11704
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51092 354 51120 11698
rect 52472 6914 52500 260102
rect 52552 229764 52604 229770
rect 52552 229706 52604 229712
rect 52564 16574 52592 229706
rect 53852 16574 53880 326334
rect 84200 319456 84252 319462
rect 84200 319398 84252 319404
rect 60740 316736 60792 316742
rect 60740 316678 60792 316684
rect 57980 313948 58032 313954
rect 57980 313890 58032 313896
rect 56600 228404 56652 228410
rect 56600 228346 56652 228352
rect 55220 36576 55272 36582
rect 55220 36518 55272 36524
rect 55232 16574 55260 36518
rect 56612 16574 56640 228346
rect 57992 16574 58020 313890
rect 59360 246356 59412 246362
rect 59360 246298 59412 246304
rect 52564 16546 53328 16574
rect 53852 16546 54984 16574
rect 55232 16546 56088 16574
rect 56612 16546 56824 16574
rect 57992 16546 58480 16574
rect 52472 6886 52592 6914
rect 52564 480 52592 6886
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53300 354 53328 16546
rect 54956 480 54984 16546
rect 56060 480 56088 16546
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58452 480 58480 16546
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 246298
rect 60752 3330 60780 316678
rect 66260 315308 66312 315314
rect 66260 315250 66312 315256
rect 60832 287700 60884 287706
rect 60832 287642 60884 287648
rect 60740 3324 60792 3330
rect 60740 3266 60792 3272
rect 60844 480 60872 287642
rect 64880 280832 64932 280838
rect 64880 280774 64932 280780
rect 63500 269816 63552 269822
rect 63500 269758 63552 269764
rect 62120 244928 62172 244934
rect 62120 244870 62172 244876
rect 62132 16574 62160 244870
rect 63512 16574 63540 269758
rect 64892 16574 64920 280774
rect 66272 16574 66300 315250
rect 77300 309800 77352 309806
rect 77300 309742 77352 309748
rect 75920 307080 75972 307086
rect 75920 307022 75972 307028
rect 70400 268388 70452 268394
rect 70400 268330 70452 268336
rect 69020 254584 69072 254590
rect 69020 254526 69072 254532
rect 67640 227044 67692 227050
rect 67640 226986 67692 226992
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 64892 16546 65104 16574
rect 66272 16546 66760 16574
rect 61660 3324 61712 3330
rect 61660 3266 61712 3272
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61672 354 61700 3266
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 61998 354 62110 480
rect 61672 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66732 480 66760 16546
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 226986
rect 69032 6914 69060 254526
rect 69112 39364 69164 39370
rect 69112 39306 69164 39312
rect 69124 16574 69152 39306
rect 70412 16574 70440 268330
rect 73160 243568 73212 243574
rect 73160 243510 73212 243516
rect 73172 16574 73200 243510
rect 74540 225616 74592 225622
rect 74540 225558 74592 225564
rect 74552 16574 74580 225558
rect 69124 16546 69888 16574
rect 70412 16546 71544 16574
rect 73172 16546 73384 16574
rect 74552 16546 75040 16574
rect 69032 6886 69152 6914
rect 69124 480 69152 6886
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 16546
rect 71516 480 71544 16546
rect 72608 10328 72660 10334
rect 72608 10270 72660 10276
rect 72620 480 72648 10270
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75012 480 75040 16546
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 307022
rect 77312 6914 77340 309742
rect 78680 284980 78732 284986
rect 78680 284922 78732 284928
rect 77392 42084 77444 42090
rect 77392 42026 77444 42032
rect 77404 16574 77432 42026
rect 78692 16574 78720 284922
rect 81440 275324 81492 275330
rect 81440 275266 81492 275272
rect 80060 242208 80112 242214
rect 80060 242150 80112 242156
rect 80072 16574 80100 242150
rect 81452 16574 81480 275266
rect 82820 253224 82872 253230
rect 82820 253166 82872 253172
rect 82832 16574 82860 253166
rect 77404 16546 78168 16574
rect 78692 16546 79272 16574
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 77312 6886 77432 6914
rect 77404 480 77432 6886
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 16546
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 319398
rect 85592 3330 85620 327694
rect 88340 304292 88392 304298
rect 88340 304234 88392 304240
rect 85672 221468 85724 221474
rect 85672 221410 85724 221416
rect 85580 3324 85632 3330
rect 85580 3266 85632 3272
rect 85684 480 85712 221410
rect 88352 16574 88380 304234
rect 89720 283620 89772 283626
rect 89720 283562 89772 283568
rect 89732 16574 89760 283562
rect 90376 202842 90404 329015
rect 93860 318096 93912 318102
rect 93860 318038 93912 318044
rect 92480 220108 92532 220114
rect 92480 220050 92532 220056
rect 90364 202836 90416 202842
rect 90364 202778 90416 202784
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 87512 15904 87564 15910
rect 87512 15846 87564 15852
rect 86500 3324 86552 3330
rect 86500 3266 86552 3272
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86512 354 86540 3266
rect 86838 354 86950 480
rect 86512 326 86950 354
rect 87524 354 87552 15846
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91560 15972 91612 15978
rect 91560 15914 91612 15920
rect 91572 480 91600 15914
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 220050
rect 93872 6914 93900 318038
rect 96620 286340 96672 286346
rect 96620 286282 96672 286288
rect 93952 239420 94004 239426
rect 93952 239362 94004 239368
rect 93964 16574 93992 239362
rect 95240 47592 95292 47598
rect 95240 47534 95292 47540
rect 95252 16574 95280 47534
rect 96632 16574 96660 286282
rect 98012 16574 98040 331842
rect 103520 330540 103572 330546
rect 103520 330482 103572 330488
rect 102140 297424 102192 297430
rect 102140 297366 102192 297372
rect 99380 273964 99432 273970
rect 99380 273906 99432 273912
rect 99392 16574 99420 273906
rect 100760 251864 100812 251870
rect 100760 251806 100812 251812
rect 93964 16546 94728 16574
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 93872 6886 93992 6914
rect 93964 480 93992 6886
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94700 354 94728 16546
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 251806
rect 102152 6914 102180 297366
rect 102232 218748 102284 218754
rect 102232 218690 102284 218696
rect 102244 16574 102272 218690
rect 103532 16574 103560 330482
rect 106280 272536 106332 272542
rect 106280 272478 106332 272484
rect 106292 16574 106320 272478
rect 102244 16546 103376 16574
rect 103532 16546 104112 16574
rect 106292 16546 106504 16574
rect 102152 6886 102272 6914
rect 102244 480 102272 6886
rect 103348 480 103376 16546
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105728 16040 105780 16046
rect 105728 15982 105780 15988
rect 105740 480 105768 15982
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 109040 16108 109092 16114
rect 109040 16050 109092 16056
rect 108120 14476 108172 14482
rect 108120 14418 108172 14424
rect 108132 480 108160 14418
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109052 354 109080 16050
rect 110432 6914 110460 336058
rect 110512 300144 110564 300150
rect 110512 300086 110564 300092
rect 110524 16574 110552 300086
rect 114560 290488 114612 290494
rect 114560 290430 114612 290436
rect 111800 238060 111852 238066
rect 111800 238002 111852 238008
rect 111812 16574 111840 238002
rect 113180 49020 113232 49026
rect 113180 48962 113232 48968
rect 113192 16574 113220 48962
rect 114572 16574 114600 290430
rect 115940 236700 115992 236706
rect 115940 236642 115992 236648
rect 115952 16574 115980 236642
rect 110524 16546 111656 16574
rect 111812 16546 112392 16574
rect 113192 16546 114048 16574
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 110432 6886 110552 6914
rect 110524 480 110552 6886
rect 111628 480 111656 16546
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114020 480 114048 16546
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 336126
rect 205640 334756 205692 334762
rect 205640 334698 205692 334704
rect 160100 334688 160152 334694
rect 160100 334630 160152 334636
rect 125600 333328 125652 333334
rect 125600 333270 125652 333276
rect 118700 250504 118752 250510
rect 118700 250446 118752 250452
rect 118712 6914 118740 250446
rect 122840 43444 122892 43450
rect 122840 43386 122892 43392
rect 118792 17264 118844 17270
rect 118792 17206 118844 17212
rect 118804 16574 118832 17206
rect 122852 16574 122880 43386
rect 118804 16546 119936 16574
rect 122852 16546 123064 16574
rect 118712 6886 118832 6914
rect 118804 480 118832 6886
rect 119908 480 119936 16546
rect 122288 14544 122340 14550
rect 122288 14486 122340 14492
rect 121092 3324 121144 3330
rect 121092 3266 121144 3272
rect 121104 480 121132 3266
rect 122300 480 122328 14486
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124680 3256 124732 3262
rect 124680 3198 124732 3204
rect 124692 480 124720 3198
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125612 354 125640 333270
rect 149060 329112 149112 329118
rect 149060 329054 149112 329060
rect 142160 322312 142212 322318
rect 142160 322254 142212 322260
rect 131120 320884 131172 320890
rect 131120 320826 131172 320832
rect 128360 315376 128412 315382
rect 128360 315318 128412 315324
rect 126980 297492 127032 297498
rect 126980 297434 127032 297440
rect 126992 480 127020 297434
rect 127072 51740 127124 51746
rect 127072 51682 127124 51688
rect 127084 16574 127112 51682
rect 128372 16574 128400 315318
rect 129740 287768 129792 287774
rect 129740 287710 129792 287716
rect 129752 16574 129780 287710
rect 131132 16574 131160 320826
rect 135260 312656 135312 312662
rect 135260 312598 135312 312604
rect 133880 282192 133932 282198
rect 133880 282134 133932 282140
rect 127084 16546 128216 16574
rect 128372 16546 128952 16574
rect 129752 16546 130608 16574
rect 131132 16546 131344 16574
rect 128188 480 128216 16546
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 130580 480 130608 16546
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 132960 8968 133012 8974
rect 132960 8910 133012 8916
rect 132972 480 133000 8910
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 133892 354 133920 282134
rect 135272 4214 135300 312598
rect 139400 305720 139452 305726
rect 139400 305662 139452 305668
rect 135352 261520 135404 261526
rect 135352 261462 135404 261468
rect 135260 4208 135312 4214
rect 135260 4150 135312 4156
rect 135364 3482 135392 261462
rect 138020 258732 138072 258738
rect 138020 258674 138072 258680
rect 138032 16574 138060 258674
rect 139412 16574 139440 305662
rect 140780 37936 140832 37942
rect 140780 37878 140832 37884
rect 140792 16574 140820 37878
rect 138032 16546 138888 16574
rect 139412 16546 139624 16574
rect 140792 16546 141280 16574
rect 137192 13116 137244 13122
rect 137192 13058 137244 13064
rect 136456 4208 136508 4214
rect 136456 4150 136508 4156
rect 135272 3454 135392 3482
rect 135272 480 135300 3454
rect 136468 480 136496 4150
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 13058
rect 138860 480 138888 16546
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 141252 480 141280 16546
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142172 354 142200 322254
rect 147680 309868 147732 309874
rect 147680 309810 147732 309816
rect 143540 308508 143592 308514
rect 143540 308450 143592 308456
rect 143552 11830 143580 308450
rect 143632 304360 143684 304366
rect 143632 304302 143684 304308
rect 143540 11824 143592 11830
rect 143540 11766 143592 11772
rect 143644 6914 143672 304302
rect 146300 303000 146352 303006
rect 146300 302942 146352 302948
rect 144920 257372 144972 257378
rect 144920 257314 144972 257320
rect 144932 16574 144960 257314
rect 146312 16574 146340 302942
rect 147692 16574 147720 309810
rect 149072 16574 149100 329054
rect 155960 323672 156012 323678
rect 155960 323614 156012 323620
rect 150440 301572 150492 301578
rect 150440 301514 150492 301520
rect 150452 16574 150480 301514
rect 153200 300212 153252 300218
rect 153200 300154 153252 300160
rect 151820 276684 151872 276690
rect 151820 276626 151872 276632
rect 144932 16546 145512 16574
rect 146312 16546 147168 16574
rect 147692 16546 147904 16574
rect 149072 16546 149560 16574
rect 150452 16546 150664 16574
rect 144736 11824 144788 11830
rect 144736 11766 144788 11772
rect 143552 6886 143672 6914
rect 143552 480 143580 6886
rect 144748 480 144776 11766
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 147140 480 147168 16546
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 149532 480 149560 16546
rect 150636 480 150664 16546
rect 151832 480 151860 276626
rect 151912 256012 151964 256018
rect 151912 255954 151964 255960
rect 151924 16574 151952 255954
rect 153212 16574 153240 300154
rect 154580 22772 154632 22778
rect 154580 22714 154632 22720
rect 154592 16574 154620 22714
rect 155972 16574 156000 323614
rect 157340 298852 157392 298858
rect 157340 298794 157392 298800
rect 157352 16574 157380 298794
rect 158720 222896 158772 222902
rect 158720 222838 158772 222844
rect 158732 16574 158760 222838
rect 151924 16546 153056 16574
rect 153212 16546 153792 16574
rect 154592 16546 155448 16574
rect 155972 16546 156184 16574
rect 157352 16546 157840 16574
rect 158732 16546 158944 16574
rect 153028 480 153056 16546
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16546
rect 155420 480 155448 16546
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 157812 480 157840 16546
rect 158916 480 158944 16546
rect 160112 11830 160140 334630
rect 189080 327888 189132 327894
rect 189080 327830 189132 327836
rect 161480 327820 161532 327826
rect 161480 327762 161532 327768
rect 160192 35216 160244 35222
rect 160192 35158 160244 35164
rect 160100 11824 160152 11830
rect 160100 11766 160152 11772
rect 160204 6914 160232 35158
rect 161492 16574 161520 327762
rect 182180 326460 182232 326466
rect 182180 326402 182232 326408
rect 164240 325032 164292 325038
rect 164240 324974 164292 324980
rect 162860 275392 162912 275398
rect 162860 275334 162912 275340
rect 162872 16574 162900 275334
rect 164252 16574 164280 324974
rect 171140 323740 171192 323746
rect 171140 323682 171192 323688
rect 165620 296064 165672 296070
rect 165620 296006 165672 296012
rect 165632 16574 165660 296006
rect 167000 274032 167052 274038
rect 167000 273974 167052 273980
rect 167012 16574 167040 273974
rect 169760 272604 169812 272610
rect 169760 272546 169812 272552
rect 169772 16574 169800 272546
rect 171152 16574 171180 323682
rect 175280 322380 175332 322386
rect 175280 322322 175332 322328
rect 173900 271176 173952 271182
rect 173900 271118 173952 271124
rect 172520 18624 172572 18630
rect 172520 18566 172572 18572
rect 172532 16574 172560 18566
rect 161492 16546 162072 16574
rect 162872 16546 163728 16574
rect 164252 16546 164464 16574
rect 165632 16546 166120 16574
rect 167012 16546 167224 16574
rect 169772 16546 170352 16574
rect 171152 16546 172008 16574
rect 172532 16546 172744 16574
rect 161296 11824 161348 11830
rect 161296 11766 161348 11772
rect 160112 6886 160232 6914
rect 160112 480 160140 6886
rect 161308 480 161336 11766
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 16546
rect 163700 480 163728 16546
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164436 354 164464 16546
rect 166092 480 166120 16546
rect 167196 480 167224 16546
rect 169576 6180 169628 6186
rect 169576 6122 169628 6128
rect 168380 4820 168432 4826
rect 168380 4762 168432 4768
rect 168392 480 168420 4762
rect 169588 480 169616 6122
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 16546
rect 171980 480 172008 16546
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173912 354 173940 271118
rect 175292 16574 175320 322322
rect 178040 320952 178092 320958
rect 178040 320894 178092 320900
rect 176660 294704 176712 294710
rect 176660 294646 176712 294652
rect 175292 16546 175504 16574
rect 175476 480 175504 16546
rect 176672 480 176700 294646
rect 176752 24132 176804 24138
rect 176752 24074 176804 24080
rect 176764 16574 176792 24074
rect 178052 16574 178080 320894
rect 179420 307148 179472 307154
rect 179420 307090 179472 307096
rect 179432 16574 179460 307090
rect 180800 269884 180852 269890
rect 180800 269826 180852 269832
rect 180812 16574 180840 269826
rect 176764 16546 177896 16574
rect 178052 16546 178632 16574
rect 179432 16546 180288 16574
rect 180812 16546 181024 16574
rect 177868 480 177896 16546
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 173134 -960 173246 326
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 180260 480 180288 16546
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 326402
rect 184940 318164 184992 318170
rect 184940 318106 184992 318112
rect 183560 291916 183612 291922
rect 183560 291858 183612 291864
rect 183572 16574 183600 291858
rect 183572 16546 183784 16574
rect 183756 480 183784 16546
rect 184952 11830 184980 318106
rect 185032 268456 185084 268462
rect 185032 268398 185084 268404
rect 184940 11824 184992 11830
rect 184940 11766 184992 11772
rect 185044 6914 185072 268398
rect 187700 265668 187752 265674
rect 187700 265610 187752 265616
rect 186320 25560 186372 25566
rect 186320 25502 186372 25508
rect 186332 16574 186360 25502
rect 187712 16574 187740 265610
rect 189092 16574 189120 327830
rect 201500 326528 201552 326534
rect 201500 326470 201552 326476
rect 200120 319524 200172 319530
rect 200120 319466 200172 319472
rect 197360 318232 197412 318238
rect 197360 318174 197412 318180
rect 193220 316804 193272 316810
rect 193220 316746 193272 316752
rect 190460 290556 190512 290562
rect 190460 290498 190512 290504
rect 186332 16546 186912 16574
rect 187712 16546 188568 16574
rect 189092 16546 189304 16574
rect 186136 11824 186188 11830
rect 186136 11766 186188 11772
rect 184952 6886 185072 6914
rect 184952 480 184980 6886
rect 186148 480 186176 11766
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 188540 480 188568 16546
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189276 354 189304 16546
rect 189694 354 189806 480
rect 189276 326 189806 354
rect 190472 354 190500 290498
rect 191840 264240 191892 264246
rect 191840 264182 191892 264188
rect 191852 16574 191880 264182
rect 191852 16546 192064 16574
rect 192036 480 192064 16546
rect 193232 480 193260 316746
rect 195980 314016 196032 314022
rect 195980 313958 196032 313964
rect 193312 289196 193364 289202
rect 193312 289138 193364 289144
rect 193324 16574 193352 289138
rect 194600 26920 194652 26926
rect 194600 26862 194652 26868
rect 194612 16574 194640 26862
rect 195992 16574 196020 313958
rect 197372 16574 197400 318174
rect 198740 262948 198792 262954
rect 198740 262890 198792 262896
rect 193324 16546 194456 16574
rect 194612 16546 195192 16574
rect 195992 16546 196848 16574
rect 197372 16546 197952 16574
rect 194428 480 194456 16546
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 189694 -960 189806 326
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 196820 480 196848 16546
rect 197924 480 197952 16546
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 262890
rect 200132 16574 200160 319466
rect 200132 16546 200344 16574
rect 200316 480 200344 16546
rect 201512 480 201540 326470
rect 202880 311228 202932 311234
rect 202880 311170 202932 311176
rect 201592 304428 201644 304434
rect 201592 304370 201644 304376
rect 201604 16574 201632 304370
rect 202892 16574 202920 311170
rect 204260 21412 204312 21418
rect 204260 21354 204312 21360
rect 204272 16574 204300 21354
rect 205652 16574 205680 334698
rect 207020 331968 207072 331974
rect 207020 331910 207072 331916
rect 201604 16546 202736 16574
rect 202892 16546 203472 16574
rect 204272 16546 205128 16574
rect 205652 16546 206232 16574
rect 202708 480 202736 16546
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 16546
rect 205100 480 205128 16546
rect 206204 480 206232 16546
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 331910
rect 213920 330608 213972 330614
rect 213920 330550 213972 330556
rect 211160 315444 211212 315450
rect 211160 315386 211212 315392
rect 209780 309936 209832 309942
rect 209780 309878 209832 309884
rect 208400 286408 208452 286414
rect 208400 286350 208452 286356
rect 208412 16574 208440 286350
rect 208412 16546 208624 16574
rect 208596 480 208624 16546
rect 209792 9674 209820 309878
rect 209872 28280 209924 28286
rect 209872 28222 209924 28228
rect 209700 9654 209820 9674
rect 209688 9648 209820 9654
rect 209740 9646 209820 9648
rect 209688 9590 209740 9596
rect 209884 6914 209912 28222
rect 211172 16574 211200 315386
rect 212540 29640 212592 29646
rect 212540 29582 212592 29588
rect 212552 16574 212580 29582
rect 213932 16574 213960 330550
rect 215300 293276 215352 293282
rect 215300 293218 215352 293224
rect 211172 16546 211752 16574
rect 212552 16546 213408 16574
rect 213932 16546 214512 16574
rect 210976 9648 211028 9654
rect 210976 9590 211028 9596
rect 209792 6886 209912 6914
rect 209792 480 209820 6886
rect 210988 480 211016 9590
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 213380 480 213408 16546
rect 214484 480 214512 16546
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 293218
rect 217336 189038 217364 463830
rect 218060 316872 218112 316878
rect 218060 316814 218112 316820
rect 217324 189032 217376 189038
rect 217324 188974 217376 188980
rect 216680 188352 216732 188358
rect 216680 188294 216732 188300
rect 216692 16574 216720 188294
rect 216692 16546 216904 16574
rect 216876 480 216904 16546
rect 218072 4214 218100 316814
rect 219440 303068 219492 303074
rect 219440 303010 219492 303016
rect 219452 16574 219480 303010
rect 220096 241466 220124 463898
rect 235356 462868 235408 462874
rect 235356 462810 235408 462816
rect 221464 462732 221516 462738
rect 221464 462674 221516 462680
rect 220820 333396 220872 333402
rect 220820 333338 220872 333344
rect 220084 241460 220136 241466
rect 220084 241402 220136 241408
rect 220832 16574 220860 333338
rect 221476 293962 221504 462674
rect 229744 461372 229796 461378
rect 229744 461314 229796 461320
rect 228364 461168 228416 461174
rect 228364 461110 228416 461116
rect 224224 461100 224276 461106
rect 224224 461042 224276 461048
rect 223580 312724 223632 312730
rect 223580 312666 223632 312672
rect 221464 293956 221516 293962
rect 221464 293898 221516 293904
rect 222200 285048 222252 285054
rect 222200 284990 222252 284996
rect 222212 16574 222240 284990
rect 219452 16546 220032 16574
rect 220832 16546 221136 16574
rect 222212 16546 222792 16574
rect 218152 7676 218204 7682
rect 218152 7618 218204 7624
rect 218060 4208 218112 4214
rect 218060 4150 218112 4156
rect 218164 3482 218192 7618
rect 219256 4208 219308 4214
rect 219256 4150 219308 4156
rect 218072 3454 218192 3482
rect 218072 480 218100 3454
rect 219268 480 219296 4150
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 16546
rect 222764 480 222792 16546
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 312666
rect 224236 33114 224264 461042
rect 225604 458380 225656 458386
rect 225604 458322 225656 458328
rect 224960 329180 225012 329186
rect 224960 329122 225012 329128
rect 224224 33108 224276 33114
rect 224224 33050 224276 33056
rect 224972 16574 225000 329122
rect 225616 71738 225644 458322
rect 227720 308576 227772 308582
rect 227720 308518 227772 308524
rect 226340 283688 226392 283694
rect 226340 283630 226392 283636
rect 225604 71732 225656 71738
rect 225604 71674 225656 71680
rect 224972 16546 225184 16574
rect 225156 480 225184 16546
rect 226352 480 226380 283630
rect 226432 31068 226484 31074
rect 226432 31010 226484 31016
rect 226444 16574 226472 31010
rect 227732 16574 227760 308518
rect 228376 111790 228404 461110
rect 229100 314084 229152 314090
rect 229100 314026 229152 314032
rect 228364 111784 228416 111790
rect 228364 111726 228416 111732
rect 229112 16574 229140 314026
rect 229756 164218 229784 461314
rect 235264 458924 235316 458930
rect 235264 458866 235316 458872
rect 233976 458720 234028 458726
rect 233976 458662 234028 458668
rect 232504 458652 232556 458658
rect 232504 458594 232556 458600
rect 231860 325100 231912 325106
rect 231860 325042 231912 325048
rect 230480 301640 230532 301646
rect 230480 301582 230532 301588
rect 229744 164212 229796 164218
rect 229744 164154 229796 164160
rect 230492 16574 230520 301582
rect 226444 16546 227576 16574
rect 227732 16546 228312 16574
rect 229112 16546 229416 16574
rect 230492 16546 231072 16574
rect 227548 480 227576 16546
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16546
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 16546
rect 231044 480 231072 16546
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 325042
rect 232516 267714 232544 458594
rect 233884 336524 233936 336530
rect 233884 336466 233936 336472
rect 233240 280900 233292 280906
rect 233240 280842 233292 280848
rect 232504 267708 232556 267714
rect 232504 267650 232556 267656
rect 233252 16574 233280 280842
rect 233252 16546 233464 16574
rect 233436 480 233464 16546
rect 233896 7614 233924 336466
rect 233988 320142 234016 458662
rect 235276 372570 235304 458866
rect 235368 411262 235396 462810
rect 264888 462800 264940 462806
rect 264888 462742 264940 462748
rect 260380 462664 260432 462670
rect 260380 462606 260432 462612
rect 247868 462528 247920 462534
rect 247868 462470 247920 462476
rect 242808 462460 242860 462466
rect 242808 462402 242860 462408
rect 236736 461440 236788 461446
rect 236736 461382 236788 461388
rect 236012 457286 236624 457314
rect 235356 411256 235408 411262
rect 235356 411198 235408 411204
rect 236012 398970 236040 457286
rect 236748 402974 236776 461382
rect 241428 458312 241480 458318
rect 241428 458254 241480 458260
rect 241440 457994 241468 458254
rect 241316 457966 241468 457994
rect 242820 457994 242848 462402
rect 246304 458448 246356 458454
rect 246304 458390 246356 458396
rect 246316 457994 246344 458390
rect 247880 457994 247908 462470
rect 250904 461304 250956 461310
rect 250904 461246 250956 461252
rect 250916 457994 250944 461246
rect 257252 461236 257304 461242
rect 257252 461178 257304 461184
rect 255688 458584 255740 458590
rect 255688 458526 255740 458532
rect 255700 457994 255728 458526
rect 257264 457994 257292 461178
rect 260392 457994 260420 462606
rect 264900 457994 264928 462742
rect 266372 460086 266400 697546
rect 298100 643136 298152 643142
rect 298100 643078 298152 643084
rect 296720 616888 296772 616894
rect 296720 616830 296772 616836
rect 293960 590708 294012 590714
rect 293960 590650 294012 590656
rect 292580 563100 292632 563106
rect 292580 563042 292632 563048
rect 288440 536852 288492 536858
rect 288440 536794 288492 536800
rect 287060 510672 287112 510678
rect 287060 510614 287112 510620
rect 284300 484424 284352 484430
rect 284300 484366 284352 484372
rect 284312 480254 284340 484366
rect 287072 480254 287100 510614
rect 288452 480254 288480 536794
rect 291200 524476 291252 524482
rect 291200 524418 291252 524424
rect 284312 480226 284708 480254
rect 287072 480226 287836 480254
rect 288452 480226 289400 480254
rect 277216 464092 277268 464098
rect 277216 464034 277268 464040
rect 269764 461032 269816 461038
rect 269764 460974 269816 460980
rect 266360 460080 266412 460086
rect 266360 460022 266412 460028
rect 266268 458516 266320 458522
rect 266268 458458 266320 458464
rect 242820 457966 242880 457994
rect 246008 457966 246344 457994
rect 247572 457966 247908 457994
rect 250700 457966 250944 457994
rect 255392 457966 255728 457994
rect 256956 457966 257292 457994
rect 260084 457966 260420 457994
rect 264776 457966 264928 457994
rect 266280 457994 266308 458458
rect 269776 457994 269804 460974
rect 274456 458788 274508 458794
rect 274456 458730 274508 458736
rect 274468 457994 274496 458730
rect 266280 457966 266340 457994
rect 269468 457966 269804 457994
rect 274160 457966 274496 457994
rect 277228 457858 277256 464034
rect 280712 463820 280764 463826
rect 280712 463762 280764 463768
rect 279148 462596 279200 462602
rect 279148 462538 279200 462544
rect 279160 457994 279188 462538
rect 280724 457994 280752 463762
rect 282276 459604 282328 459610
rect 282276 459546 282328 459552
rect 282288 457994 282316 459546
rect 278852 457966 279188 457994
rect 280416 457966 280752 457994
rect 281980 457966 282316 457994
rect 284680 457994 284708 480226
rect 286232 470620 286284 470626
rect 286232 470562 286284 470568
rect 286244 457994 286272 470562
rect 287808 457994 287836 480226
rect 289372 457994 289400 480226
rect 291212 457994 291240 524418
rect 292592 457994 292620 563042
rect 293972 480254 294000 590650
rect 295340 576904 295392 576910
rect 295340 576846 295392 576852
rect 295352 480254 295380 576846
rect 296732 480254 296760 616830
rect 298112 480254 298140 643078
rect 299480 630692 299532 630698
rect 299480 630634 299532 630640
rect 299492 480254 299520 630634
rect 293972 480226 294092 480254
rect 295352 480226 295656 480254
rect 296732 480226 297220 480254
rect 298112 480226 298784 480254
rect 299492 480226 300348 480254
rect 294064 457994 294092 480226
rect 295628 457994 295656 480226
rect 297192 457994 297220 480226
rect 298756 457994 298784 480226
rect 300320 457994 300348 480226
rect 301516 465730 301544 699994
rect 303620 696992 303672 696998
rect 303620 696934 303672 696940
rect 302240 670812 302292 670818
rect 302240 670754 302292 670760
rect 301504 465724 301556 465730
rect 301504 465666 301556 465672
rect 302252 457994 302280 670754
rect 303632 457994 303660 696934
rect 305000 683188 305052 683194
rect 305000 683130 305052 683136
rect 305012 457994 305040 683130
rect 318812 480254 318840 700606
rect 320180 502988 320232 502994
rect 320180 502930 320232 502936
rect 320192 480254 320220 502930
rect 322952 480254 322980 700742
rect 328460 700732 328512 700738
rect 328460 700674 328512 700680
rect 318812 480226 319116 480254
rect 320192 480226 320680 480254
rect 322952 480226 323808 480254
rect 311256 472660 311308 472666
rect 311256 472602 311308 472608
rect 307300 461644 307352 461650
rect 307300 461586 307352 461592
rect 307312 457994 307340 461586
rect 308864 460624 308916 460630
rect 308864 460566 308916 460572
rect 308496 459604 308548 459610
rect 308496 459546 308548 459552
rect 308508 458862 308536 459546
rect 308496 458856 308548 458862
rect 308496 458798 308548 458804
rect 308876 457994 308904 460566
rect 310428 460556 310480 460562
rect 310428 460498 310480 460504
rect 310440 457994 310468 460498
rect 284680 457966 285108 457994
rect 286244 457966 286672 457994
rect 287808 457966 288236 457994
rect 289372 457966 289800 457994
rect 291212 457966 291364 457994
rect 292592 457966 292928 457994
rect 294064 457966 294492 457994
rect 295628 457966 296056 457994
rect 297192 457966 297620 457994
rect 298756 457966 299184 457994
rect 300320 457966 300748 457994
rect 302252 457966 302312 457994
rect 303632 457966 303876 457994
rect 305012 457966 305440 457994
rect 307004 457966 307340 457994
rect 308568 457966 308904 457994
rect 310132 457966 310468 457994
rect 311268 457994 311296 472602
rect 316040 464364 316092 464370
rect 316040 464306 316092 464312
rect 313188 460828 313240 460834
rect 313188 460770 313240 460776
rect 313200 457994 313228 460770
rect 315120 460760 315172 460766
rect 315120 460702 315172 460708
rect 315132 457994 315160 460702
rect 311268 457966 311696 457994
rect 313200 457966 313260 457994
rect 314824 457966 315160 457994
rect 316052 457994 316080 464306
rect 318248 460148 318300 460154
rect 318248 460090 318300 460096
rect 318260 457994 318288 460090
rect 316052 457966 316388 457994
rect 317952 457966 318288 457994
rect 319088 457994 319116 480226
rect 320652 457994 320680 480226
rect 322848 460012 322900 460018
rect 322848 459954 322900 459960
rect 322860 457994 322888 459954
rect 319088 457966 319516 457994
rect 320652 457966 321080 457994
rect 322644 457966 322888 457994
rect 323780 457994 323808 480226
rect 325700 465724 325752 465730
rect 325700 465666 325752 465672
rect 325712 457994 325740 465666
rect 327080 460080 327132 460086
rect 327080 460022 327132 460028
rect 327092 457994 327120 460022
rect 328472 457994 328500 700674
rect 330024 467152 330076 467158
rect 330024 467094 330076 467100
rect 330036 457994 330064 467094
rect 331232 460018 331260 702986
rect 348804 700806 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 348792 700800 348844 700806
rect 348792 700742 348844 700748
rect 332600 700596 332652 700602
rect 332600 700538 332652 700544
rect 332612 480254 332640 700538
rect 338120 700528 338172 700534
rect 338120 700470 338172 700476
rect 332612 480226 333192 480254
rect 331680 460896 331732 460902
rect 331680 460838 331732 460844
rect 331220 460012 331272 460018
rect 331220 459954 331272 459960
rect 331692 457994 331720 460838
rect 333164 457994 333192 480226
rect 334716 468512 334768 468518
rect 334716 468454 334768 468460
rect 334728 457994 334756 468454
rect 336372 460692 336424 460698
rect 336372 460634 336424 460640
rect 336384 457994 336412 460634
rect 338132 457994 338160 700470
rect 342260 700460 342312 700466
rect 342260 700402 342312 700408
rect 342272 480254 342300 700402
rect 346400 700392 346452 700398
rect 346400 700334 346452 700340
rect 345020 700324 345072 700330
rect 345020 700266 345072 700272
rect 345032 480254 345060 700266
rect 346412 480254 346440 700334
rect 351920 670744 351972 670750
rect 351920 670686 351972 670692
rect 350540 656940 350592 656946
rect 350540 656882 350592 656888
rect 342272 480226 342576 480254
rect 345032 480226 345704 480254
rect 346412 480226 347268 480254
rect 339500 469872 339552 469878
rect 339500 469814 339552 469820
rect 339512 457994 339540 469814
rect 341064 460488 341116 460494
rect 341064 460430 341116 460436
rect 341076 457994 341104 460430
rect 342548 457994 342576 480226
rect 344100 474020 344152 474026
rect 344100 473962 344152 473968
rect 344112 457994 344140 473962
rect 345676 457994 345704 480226
rect 347240 457994 347268 480226
rect 349158 460184 349214 460193
rect 349158 460119 349214 460128
rect 349172 457994 349200 460119
rect 350552 457994 350580 656882
rect 351932 457994 351960 670686
rect 356060 618316 356112 618322
rect 356060 618258 356112 618264
rect 354680 605872 354732 605878
rect 354680 605814 354732 605820
rect 354692 480254 354720 605814
rect 356072 480254 356100 618258
rect 361580 565888 361632 565894
rect 361580 565830 361632 565836
rect 358820 553444 358872 553450
rect 358820 553386 358872 553392
rect 358832 480254 358860 553386
rect 354692 480226 355088 480254
rect 356072 480226 356652 480254
rect 358832 480226 359780 480254
rect 353576 460420 353628 460426
rect 353576 460362 353628 460368
rect 353300 459604 353352 459610
rect 353300 459546 353352 459552
rect 323780 457966 324208 457994
rect 325712 457966 325772 457994
rect 327092 457966 327336 457994
rect 328472 457966 328900 457994
rect 330036 457966 330464 457994
rect 331692 457966 332028 457994
rect 333164 457966 333592 457994
rect 334728 457966 335156 457994
rect 336384 457966 336720 457994
rect 338132 457966 338284 457994
rect 339512 457966 339848 457994
rect 341076 457966 341412 457994
rect 342548 457966 342976 457994
rect 344112 457966 344540 457994
rect 345676 457966 346104 457994
rect 347240 457966 347668 457994
rect 349172 457966 349232 457994
rect 350552 457966 350796 457994
rect 351932 457966 352360 457994
rect 277228 457830 277288 457858
rect 235828 398942 236040 398970
rect 236104 402946 236776 402974
rect 237392 457694 238188 457722
rect 235828 398698 235856 398942
rect 236104 398834 236132 402946
rect 235920 398818 236132 398834
rect 235908 398812 236132 398818
rect 235960 398806 236132 398812
rect 235908 398754 235960 398760
rect 235828 398670 236040 398698
rect 235264 372564 235316 372570
rect 235264 372506 235316 372512
rect 234620 334824 234672 334830
rect 234620 334766 234672 334772
rect 233976 320136 234028 320142
rect 233976 320078 234028 320084
rect 234632 11830 234660 334766
rect 234712 267028 234764 267034
rect 234712 266970 234764 266976
rect 234620 11824 234672 11830
rect 234620 11766 234672 11772
rect 233884 7608 233936 7614
rect 233884 7550 233936 7556
rect 234724 6914 234752 266970
rect 235816 11824 235868 11830
rect 235816 11766 235868 11772
rect 234632 6886 234752 6914
rect 234632 480 234660 6886
rect 235828 480 235856 11766
rect 236012 6866 236040 398670
rect 236092 311296 236144 311302
rect 236092 311238 236144 311244
rect 236104 16574 236132 311238
rect 237392 33114 237420 457694
rect 239416 457570 239752 457586
rect 238024 457564 238076 457570
rect 238024 457506 238076 457512
rect 239404 457564 239752 457570
rect 239456 457558 239752 457564
rect 239404 457506 239456 457512
rect 237472 240780 237524 240786
rect 237472 240722 237524 240728
rect 237380 33108 237432 33114
rect 237380 33050 237432 33056
rect 237484 16574 237512 240722
rect 238036 46238 238064 457506
rect 353312 457502 353340 459546
rect 353588 457994 353616 460362
rect 355060 457994 355088 480226
rect 356624 457994 356652 480226
rect 358268 460352 358320 460358
rect 358268 460294 358320 460300
rect 358280 457994 358308 460294
rect 359752 457994 359780 480226
rect 361592 457994 361620 565830
rect 364352 502994 364380 702406
rect 365720 514820 365772 514826
rect 365720 514762 365772 514768
rect 364340 502988 364392 502994
rect 364340 502930 364392 502936
rect 364340 501016 364392 501022
rect 364340 500958 364392 500964
rect 364352 480254 364380 500958
rect 365732 480254 365760 514762
rect 364352 480226 364472 480254
rect 365732 480226 366036 480254
rect 362960 460284 363012 460290
rect 362960 460226 363012 460232
rect 362972 457994 363000 460226
rect 364444 457994 364472 480226
rect 366008 457994 366036 480226
rect 380072 464024 380124 464030
rect 380072 463966 380124 463972
rect 378508 463752 378560 463758
rect 378508 463694 378560 463700
rect 375472 462868 375524 462874
rect 375472 462810 375524 462816
rect 370780 462392 370832 462398
rect 370780 462334 370832 462340
rect 367652 460216 367704 460222
rect 367652 460158 367704 460164
rect 367664 457994 367692 460158
rect 369216 459604 369268 459610
rect 369216 459546 369268 459552
rect 369228 457994 369256 459546
rect 370792 457994 370820 462334
rect 374000 461440 374052 461446
rect 374000 461382 374052 461388
rect 372666 458244 372718 458250
rect 372666 458186 372718 458192
rect 353588 457966 353924 457994
rect 355060 457966 355488 457994
rect 356624 457966 357052 457994
rect 358280 457966 358616 457994
rect 359752 457966 360180 457994
rect 361592 457966 361744 457994
rect 362972 457966 363308 457994
rect 364444 457966 364872 457994
rect 366008 457966 366436 457994
rect 367664 457966 368000 457994
rect 369228 457966 369564 457994
rect 370792 457966 371128 457994
rect 372678 457980 372706 458186
rect 374012 457994 374040 461382
rect 375484 457994 375512 462810
rect 377036 458924 377088 458930
rect 377036 458866 377088 458872
rect 377048 457994 377076 458866
rect 378520 457994 378548 463694
rect 380084 457994 380112 463966
rect 387892 463956 387944 463962
rect 387892 463898 387944 463904
rect 383292 462732 383344 462738
rect 383292 462674 383344 462680
rect 381728 458720 381780 458726
rect 381728 458662 381780 458668
rect 381740 457994 381768 458662
rect 383304 457994 383332 462674
rect 386420 458652 386472 458658
rect 386420 458594 386472 458600
rect 386432 457994 386460 458594
rect 387904 457994 387932 463898
rect 392584 463888 392636 463894
rect 392584 463830 392636 463836
rect 391112 460964 391164 460970
rect 391112 460906 391164 460912
rect 391124 457994 391152 460906
rect 392596 457994 392624 463830
rect 396080 461372 396132 461378
rect 396080 461314 396132 461320
rect 396092 457994 396120 461314
rect 397472 460154 397500 703520
rect 413664 700670 413692 703520
rect 413652 700664 413704 700670
rect 413652 700606 413704 700612
rect 413284 700324 413336 700330
rect 413284 700266 413336 700272
rect 413296 461650 413324 700266
rect 429856 699718 429884 703520
rect 428464 699712 428516 699718
rect 428464 699654 428516 699660
rect 429844 699712 429896 699718
rect 429844 699654 429896 699660
rect 428476 464370 428504 699654
rect 428464 464364 428516 464370
rect 428464 464306 428516 464312
rect 435364 464092 435416 464098
rect 435364 464034 435416 464040
rect 422944 462800 422996 462806
rect 422944 462742 422996 462748
rect 421564 462664 421616 462670
rect 421564 462606 421616 462612
rect 413284 461644 413336 461650
rect 413284 461586 413336 461592
rect 417424 461304 417476 461310
rect 417424 461246 417476 461252
rect 400496 461168 400548 461174
rect 400496 461110 400548 461116
rect 397460 460148 397512 460154
rect 397460 460090 397512 460096
rect 400508 457994 400536 461110
rect 409880 461100 409932 461106
rect 409880 461042 409932 461048
rect 405188 458380 405240 458386
rect 405188 458322 405240 458328
rect 405200 457994 405228 458322
rect 409892 457994 409920 461042
rect 416044 458788 416096 458794
rect 416044 458730 416096 458736
rect 414664 458448 414716 458454
rect 414664 458390 414716 458396
rect 374012 457966 374256 457994
rect 375484 457966 375820 457994
rect 377048 457966 377384 457994
rect 378520 457966 378948 457994
rect 380084 457966 380512 457994
rect 381740 457966 382076 457994
rect 383304 457966 383640 457994
rect 386432 457966 386768 457994
rect 387904 457966 388332 457994
rect 391124 457966 391460 457994
rect 392596 457966 393024 457994
rect 396092 457966 396152 457994
rect 400508 457966 400844 457994
rect 405200 457966 405536 457994
rect 409892 457966 410228 457994
rect 275928 457496 275980 457502
rect 244738 457464 244794 457473
rect 244444 457422 244738 457450
rect 244738 457399 244794 457408
rect 248970 457464 249026 457473
rect 252374 457464 252430 457473
rect 249026 457422 249136 457450
rect 252264 457422 252374 457450
rect 248970 457399 249026 457408
rect 252374 457399 252430 457408
rect 253662 457464 253718 457473
rect 258814 457464 258870 457473
rect 253718 457422 253828 457450
rect 258520 457422 258814 457450
rect 253662 457399 253718 457408
rect 261942 457464 261998 457473
rect 261648 457422 261942 457450
rect 258814 457399 258870 457408
rect 263322 457464 263378 457473
rect 263212 457422 263322 457450
rect 261942 457399 261998 457408
rect 268198 457464 268254 457473
rect 267904 457422 268198 457450
rect 263322 457399 263378 457408
rect 271326 457464 271382 457473
rect 271032 457422 271326 457450
rect 268198 457399 268254 457408
rect 272890 457464 272946 457473
rect 272596 457422 272890 457450
rect 271326 457399 271382 457408
rect 275724 457444 275928 457450
rect 283656 457496 283708 457502
rect 275724 457438 275980 457444
rect 283544 457444 283656 457450
rect 283544 457438 283708 457444
rect 353300 457496 353352 457502
rect 412088 457496 412140 457502
rect 385314 457464 385370 457473
rect 353300 457438 353352 457444
rect 275724 457422 275968 457438
rect 283544 457422 283696 457438
rect 385204 457422 385314 457450
rect 272890 457399 272946 457408
rect 385314 457399 385370 457408
rect 389638 457464 389694 457473
rect 394238 457464 394294 457473
rect 389694 457422 389896 457450
rect 389638 457399 389694 457408
rect 397550 457464 397606 457473
rect 394294 457422 394588 457450
rect 394238 457399 394294 457408
rect 398930 457464 398986 457473
rect 397606 457422 397716 457450
rect 397550 457399 397606 457408
rect 402058 457464 402114 457473
rect 398986 457422 399280 457450
rect 398930 457399 398986 457408
rect 403622 457464 403678 457473
rect 402114 457422 402408 457450
rect 402058 457399 402114 457408
rect 406750 457464 406806 457473
rect 403678 457422 403972 457450
rect 403622 457399 403678 457408
rect 408774 457464 408830 457473
rect 406806 457422 407100 457450
rect 408664 457422 408774 457450
rect 406750 457399 406806 457408
rect 411792 457444 412088 457450
rect 414112 457496 414164 457502
rect 411792 457438 412140 457444
rect 411792 457422 412128 457438
rect 413356 457422 413508 457450
rect 414112 457438 414164 457444
rect 408774 457399 408830 457408
rect 413480 451274 413508 457422
rect 413388 451246 413508 451274
rect 246302 338056 246358 338065
rect 400862 338056 400918 338065
rect 246302 337991 246358 338000
rect 256896 338014 257140 338042
rect 257264 338014 257416 338042
rect 257540 338014 257692 338042
rect 257816 338014 257968 338042
rect 243544 336388 243596 336394
rect 243544 336330 243596 336336
rect 242164 336320 242216 336326
rect 242164 336262 242216 336268
rect 238760 323808 238812 323814
rect 238760 323750 238812 323756
rect 238024 46232 238076 46238
rect 238024 46174 238076 46180
rect 238772 16574 238800 323750
rect 240140 279540 240192 279546
rect 240140 279482 240192 279488
rect 236104 16546 236592 16574
rect 237484 16546 237696 16574
rect 238772 16546 239352 16574
rect 236000 6860 236052 6866
rect 236000 6802 236052 6808
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 16546
rect 239324 480 239352 16546
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240152 354 240180 279482
rect 241520 260228 241572 260234
rect 241520 260170 241572 260176
rect 241532 16574 241560 260170
rect 241532 16546 241744 16574
rect 241716 480 241744 16546
rect 242176 6186 242204 336262
rect 242900 332036 242952 332042
rect 242900 331978 242952 331984
rect 242912 11830 242940 331978
rect 242992 322448 243044 322454
rect 242992 322390 243044 322396
rect 242900 11824 242952 11830
rect 242900 11766 242952 11772
rect 243004 6914 243032 322390
rect 243556 8974 243584 336330
rect 245660 307216 245712 307222
rect 245660 307158 245712 307164
rect 244280 33788 244332 33794
rect 244280 33730 244332 33736
rect 244292 16574 244320 33730
rect 245672 16574 245700 307158
rect 246316 60722 246344 337991
rect 256056 336728 256108 336734
rect 256056 336670 256108 336676
rect 255964 336456 256016 336462
rect 255964 336398 256016 336404
rect 247684 336252 247736 336258
rect 247684 336194 247736 336200
rect 247040 305788 247092 305794
rect 247040 305730 247092 305736
rect 246304 60716 246356 60722
rect 246304 60658 246356 60664
rect 247052 16574 247080 305730
rect 244292 16546 245240 16574
rect 245672 16546 245976 16574
rect 247052 16546 247632 16574
rect 244096 11824 244148 11830
rect 244096 11766 244148 11772
rect 243544 8968 243596 8974
rect 243544 8910 243596 8916
rect 242912 6886 243032 6914
rect 242164 6180 242216 6186
rect 242164 6122 242216 6128
rect 242912 480 242940 6886
rect 244108 480 244136 11766
rect 245212 480 245240 16546
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 16546
rect 247604 480 247632 16546
rect 247696 7682 247724 336194
rect 250442 334112 250498 334121
rect 250442 334047 250498 334056
rect 248420 333464 248472 333470
rect 248420 333406 248472 333412
rect 247684 7676 247736 7682
rect 247684 7618 247736 7624
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248432 354 248460 333406
rect 249800 321020 249852 321026
rect 249800 320962 249852 320968
rect 249812 16574 249840 320962
rect 250456 100706 250484 334047
rect 253940 330676 253992 330682
rect 253940 330618 253992 330624
rect 252560 319592 252612 319598
rect 252560 319534 252612 319540
rect 251180 278112 251232 278118
rect 251180 278054 251232 278060
rect 250444 100700 250496 100706
rect 250444 100642 250496 100648
rect 249812 16546 250024 16574
rect 249996 480 250024 16546
rect 251192 480 251220 278054
rect 251272 166320 251324 166326
rect 251272 166262 251324 166268
rect 251284 16574 251312 166262
rect 252572 16574 252600 319534
rect 253952 16574 253980 330618
rect 255320 297560 255372 297566
rect 255320 297502 255372 297508
rect 255332 16574 255360 297502
rect 251284 16546 252416 16574
rect 252572 16546 253520 16574
rect 253952 16546 254256 16574
rect 255332 16546 255912 16574
rect 252388 480 252416 16546
rect 253492 480 253520 16546
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 255884 480 255912 16546
rect 255976 4826 256004 336398
rect 256068 249082 256096 336670
rect 256148 336660 256200 336666
rect 256148 336602 256200 336608
rect 256160 289134 256188 336602
rect 256792 326392 256844 326398
rect 256792 326334 256844 326340
rect 256148 289128 256200 289134
rect 256148 289070 256200 289076
rect 256804 279478 256832 326334
rect 256896 311166 256924 338014
rect 257264 316034 257292 338014
rect 257344 336592 257396 336598
rect 257344 336534 257396 336540
rect 256988 316006 257292 316034
rect 256884 311160 256936 311166
rect 256884 311102 256936 311108
rect 256792 279472 256844 279478
rect 256792 279414 256844 279420
rect 256988 278050 257016 316006
rect 256976 278044 257028 278050
rect 256976 277986 257028 277992
rect 256056 249076 256108 249082
rect 256056 249018 256108 249024
rect 257356 11762 257384 336534
rect 257436 335368 257488 335374
rect 257436 335310 257488 335316
rect 257448 40730 257476 335310
rect 257540 326398 257568 338014
rect 257816 336734 257844 338014
rect 258230 337770 258258 338028
rect 258368 338014 258520 338042
rect 258644 338014 258796 338042
rect 258920 338014 259072 338042
rect 259196 338014 259348 338042
rect 259624 338014 259776 338042
rect 258230 337742 258304 337770
rect 257804 336728 257856 336734
rect 257804 336670 257856 336676
rect 257528 326392 257580 326398
rect 257528 326334 257580 326340
rect 258172 326392 258224 326398
rect 258172 326334 258224 326340
rect 258184 308446 258212 326334
rect 258172 308440 258224 308446
rect 258172 308382 258224 308388
rect 257436 40724 257488 40730
rect 257436 40666 257488 40672
rect 257344 11756 257396 11762
rect 257344 11698 257396 11704
rect 258276 6914 258304 337742
rect 258368 335986 258396 338014
rect 258356 335980 258408 335986
rect 258356 335922 258408 335928
rect 258644 333198 258672 338014
rect 258632 333192 258684 333198
rect 258632 333134 258684 333140
rect 258920 326398 258948 338014
rect 259196 335374 259224 338014
rect 259184 335368 259236 335374
rect 259184 335310 259236 335316
rect 258908 326392 258960 326398
rect 258908 326334 258960 326340
rect 259644 326392 259696 326398
rect 259644 326334 259696 326340
rect 259552 326256 259604 326262
rect 259552 326198 259604 326204
rect 259564 6914 259592 326198
rect 259656 224262 259684 326334
rect 259748 323626 259776 338014
rect 259840 338014 259900 338042
rect 260024 338014 260176 338042
rect 260300 338014 260452 338042
rect 260576 338014 260728 338042
rect 260852 338014 261004 338042
rect 261128 338014 261280 338042
rect 261404 338014 261556 338042
rect 261680 338014 261832 338042
rect 261956 338014 262108 338042
rect 262384 338014 262536 338042
rect 259840 334626 259868 338014
rect 260024 335354 260052 338014
rect 259932 335326 260052 335354
rect 259828 334620 259880 334626
rect 259828 334562 259880 334568
rect 259748 323598 259868 323626
rect 259736 321360 259788 321366
rect 259736 321302 259788 321308
rect 259748 301510 259776 321302
rect 259736 301504 259788 301510
rect 259736 301446 259788 301452
rect 259644 224256 259696 224262
rect 259644 224198 259696 224204
rect 259644 17332 259696 17338
rect 259644 17274 259696 17280
rect 258184 6886 258304 6914
rect 259472 6886 259592 6914
rect 255964 4820 256016 4826
rect 255964 4762 256016 4768
rect 257068 4820 257120 4826
rect 257068 4762 257120 4768
rect 257080 480 257108 4762
rect 258080 3732 258132 3738
rect 258080 3674 258132 3680
rect 258092 3194 258120 3674
rect 258184 3369 258212 6886
rect 258264 6180 258316 6186
rect 258264 6122 258316 6128
rect 258170 3360 258226 3369
rect 258170 3295 258226 3304
rect 258080 3188 258132 3194
rect 258080 3130 258132 3136
rect 258276 480 258304 6122
rect 258448 4208 258500 4214
rect 258448 4150 258500 4156
rect 258460 3602 258488 4150
rect 259472 3618 259500 6886
rect 258448 3596 258500 3602
rect 258448 3538 258500 3544
rect 259380 3590 259500 3618
rect 259380 3534 259408 3590
rect 259368 3528 259420 3534
rect 259656 3482 259684 17274
rect 259368 3470 259420 3476
rect 259472 3454 259684 3482
rect 259840 3466 259868 323598
rect 259932 321366 259960 335326
rect 260300 326398 260328 338014
rect 260288 326392 260340 326398
rect 260288 326334 260340 326340
rect 260576 326262 260604 338014
rect 260852 336666 260880 338014
rect 260840 336660 260892 336666
rect 260840 336602 260892 336608
rect 261128 335354 261156 338014
rect 261036 335326 261156 335354
rect 260564 326256 260616 326262
rect 260564 326198 260616 326204
rect 260932 326256 260984 326262
rect 260932 326198 260984 326204
rect 259920 321360 259972 321366
rect 259920 321302 259972 321308
rect 260656 7744 260708 7750
rect 260656 7686 260708 7692
rect 259828 3460 259880 3466
rect 259472 480 259500 3454
rect 259828 3402 259880 3408
rect 260668 480 260696 7686
rect 260944 3670 260972 326198
rect 261036 214606 261064 335326
rect 261208 326392 261260 326398
rect 261208 326334 261260 326340
rect 261116 324556 261168 324562
rect 261116 324498 261168 324504
rect 261128 294642 261156 324498
rect 261116 294636 261168 294642
rect 261116 294578 261168 294584
rect 261024 214600 261076 214606
rect 261024 214542 261076 214548
rect 261220 3738 261248 326334
rect 261404 326262 261432 338014
rect 261484 335708 261536 335714
rect 261484 335650 261536 335656
rect 261392 326256 261444 326262
rect 261392 326198 261444 326204
rect 261496 298790 261524 335650
rect 261680 326398 261708 338014
rect 261668 326392 261720 326398
rect 261668 326334 261720 326340
rect 261956 324562 261984 338014
rect 262312 326392 262364 326398
rect 262312 326334 262364 326340
rect 261944 324556 261996 324562
rect 261944 324498 261996 324504
rect 261484 298784 261536 298790
rect 261484 298726 261536 298732
rect 261760 9104 261812 9110
rect 261760 9046 261812 9052
rect 261208 3732 261260 3738
rect 261208 3674 261260 3680
rect 260932 3664 260984 3670
rect 260932 3606 260984 3612
rect 261772 480 261800 9046
rect 262324 3806 262352 326334
rect 262404 326256 262456 326262
rect 262404 326198 262456 326204
rect 262416 302938 262444 326198
rect 262508 323610 262536 338014
rect 262600 338014 262660 338042
rect 262784 338014 262936 338042
rect 263060 338014 263212 338042
rect 263336 338014 263488 338042
rect 263704 338014 263764 338042
rect 263888 338014 264040 338042
rect 264164 338014 264316 338042
rect 264440 338014 264592 338042
rect 264716 338014 264868 338042
rect 265144 338014 265296 338042
rect 262496 323604 262548 323610
rect 262496 323546 262548 323552
rect 262404 302932 262456 302938
rect 262404 302874 262456 302880
rect 262312 3800 262364 3806
rect 262312 3742 262364 3748
rect 262600 3194 262628 338014
rect 262784 326398 262812 338014
rect 263060 335714 263088 338014
rect 263048 335708 263100 335714
rect 263048 335650 263100 335656
rect 262772 326392 262824 326398
rect 262772 326334 262824 326340
rect 263336 326262 263364 338014
rect 263324 326256 263376 326262
rect 263324 326198 263376 326204
rect 262956 6248 263008 6254
rect 262956 6190 263008 6196
rect 262588 3188 262640 3194
rect 262588 3130 262640 3136
rect 262968 480 262996 6190
rect 263704 3874 263732 338014
rect 263888 335354 263916 338014
rect 263796 335326 263916 335354
rect 263796 326602 263824 335326
rect 264164 331214 264192 338014
rect 264244 336728 264296 336734
rect 264244 336670 264296 336676
rect 263980 331186 264192 331214
rect 263784 326596 263836 326602
rect 263784 326538 263836 326544
rect 263980 326346 264008 331186
rect 264060 326596 264112 326602
rect 264060 326538 264112 326544
rect 263796 326318 264008 326346
rect 263796 235278 263824 326318
rect 263968 326256 264020 326262
rect 263968 326198 264020 326204
rect 263876 316736 263928 316742
rect 263876 316678 263928 316684
rect 263888 291854 263916 316678
rect 263876 291848 263928 291854
rect 263876 291790 263928 291796
rect 263784 235272 263836 235278
rect 263784 235214 263836 235220
rect 263980 3942 264008 326198
rect 264072 316742 264100 326538
rect 264060 316736 264112 316742
rect 264060 316678 264112 316684
rect 264256 305658 264284 336670
rect 264440 326262 264468 338014
rect 264716 336530 264744 338014
rect 264704 336524 264756 336530
rect 264704 336466 264756 336472
rect 265268 335354 265296 338014
rect 265406 337770 265434 338028
rect 265544 338014 265696 338042
rect 265820 338014 265972 338042
rect 266096 338014 266248 338042
rect 266372 338014 266524 338042
rect 266648 338014 266800 338042
rect 266924 338014 267076 338042
rect 267200 338014 267352 338042
rect 267476 338014 267628 338042
rect 265406 337742 265480 337770
rect 265268 335326 265388 335354
rect 264980 326392 265032 326398
rect 264980 326334 265032 326340
rect 264428 326256 264480 326262
rect 264428 326198 264480 326204
rect 264244 305652 264296 305658
rect 264244 305594 264296 305600
rect 264152 8968 264204 8974
rect 264152 8910 264204 8916
rect 263968 3936 264020 3942
rect 263968 3878 264020 3884
rect 263692 3868 263744 3874
rect 263692 3810 263744 3816
rect 264164 480 264192 8910
rect 264992 4010 265020 326334
rect 265164 326256 265216 326262
rect 265164 326198 265216 326204
rect 265072 326188 265124 326194
rect 265072 326130 265124 326136
rect 265084 4078 265112 326130
rect 265176 233918 265204 326198
rect 265360 322250 265388 335326
rect 265452 326398 265480 337742
rect 265440 326392 265492 326398
rect 265440 326334 265492 326340
rect 265348 322244 265400 322250
rect 265348 322186 265400 322192
rect 265544 311894 265572 338014
rect 265820 326262 265848 338014
rect 265808 326256 265860 326262
rect 265808 326198 265860 326204
rect 266096 326194 266124 338014
rect 266372 336734 266400 338014
rect 266360 336728 266412 336734
rect 266360 336670 266412 336676
rect 266648 335354 266676 338014
rect 266556 335326 266676 335354
rect 266452 326392 266504 326398
rect 266452 326334 266504 326340
rect 266084 326188 266136 326194
rect 266084 326130 266136 326136
rect 265268 311866 265572 311894
rect 265268 296002 265296 311866
rect 265256 295996 265308 296002
rect 265256 295938 265308 295944
rect 265164 233912 265216 233918
rect 265164 233854 265216 233860
rect 266464 232558 266492 326334
rect 266556 262886 266584 335326
rect 266636 325372 266688 325378
rect 266636 325314 266688 325320
rect 266648 312594 266676 325314
rect 266636 312588 266688 312594
rect 266636 312530 266688 312536
rect 266924 311894 266952 338014
rect 267200 325378 267228 338014
rect 267476 326398 267504 338014
rect 267890 337770 267918 338028
rect 268028 338014 268180 338042
rect 268304 338014 268456 338042
rect 268580 338014 268732 338042
rect 268856 338014 269008 338042
rect 269284 338014 269436 338042
rect 267890 337742 267964 337770
rect 267464 326392 267516 326398
rect 267464 326334 267516 326340
rect 267832 326392 267884 326398
rect 267832 326334 267884 326340
rect 267936 326346 267964 337742
rect 268028 331214 268056 338014
rect 268028 331186 268148 331214
rect 267188 325372 267240 325378
rect 267188 325314 267240 325320
rect 266740 311866 266952 311894
rect 266544 262880 266596 262886
rect 266544 262822 266596 262828
rect 266452 232552 266504 232558
rect 266452 232494 266504 232500
rect 265164 11756 265216 11762
rect 265164 11698 265216 11704
rect 265072 4072 265124 4078
rect 265072 4014 265124 4020
rect 264980 4004 265032 4010
rect 264980 3946 265032 3952
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265176 354 265204 11698
rect 266544 9036 266596 9042
rect 266544 8978 266596 8984
rect 266556 480 266584 8978
rect 266740 3602 266768 311866
rect 267844 231130 267872 326334
rect 267936 326318 268056 326346
rect 267924 326256 267976 326262
rect 267924 326198 267976 326204
rect 267936 247722 267964 326198
rect 268028 321554 268056 326318
rect 268120 324970 268148 331186
rect 268304 326262 268332 338014
rect 268384 336660 268436 336666
rect 268384 336602 268436 336608
rect 268292 326256 268344 326262
rect 268292 326198 268344 326204
rect 268108 324964 268160 324970
rect 268108 324906 268160 324912
rect 268028 321526 268148 321554
rect 267924 247716 267976 247722
rect 267924 247658 267976 247664
rect 267832 231124 267884 231130
rect 267832 231066 267884 231072
rect 267740 5024 267792 5030
rect 267740 4966 267792 4972
rect 266728 3596 266780 3602
rect 266728 3538 266780 3544
rect 267752 480 267780 4966
rect 268120 3398 268148 321526
rect 268396 280838 268424 336602
rect 268580 326398 268608 338014
rect 268856 336598 268884 338014
rect 268844 336592 268896 336598
rect 268844 336534 268896 336540
rect 269408 326738 269436 338014
rect 269500 338014 269560 338042
rect 269684 338014 269836 338042
rect 269960 338014 270112 338042
rect 270236 338014 270388 338042
rect 270512 338014 270664 338042
rect 270788 338014 270940 338042
rect 271064 338014 271216 338042
rect 271340 338014 271492 338042
rect 271616 338014 271768 338042
rect 271984 338014 272044 338042
rect 272168 338014 272320 338042
rect 272444 338014 272596 338042
rect 272720 338014 272872 338042
rect 272996 338014 273148 338042
rect 273272 338014 273424 338042
rect 273548 338014 273700 338042
rect 273824 338014 273976 338042
rect 274100 338014 274252 338042
rect 274376 338014 274528 338042
rect 274804 338014 274956 338042
rect 269396 326732 269448 326738
rect 269396 326674 269448 326680
rect 269500 326602 269528 338014
rect 269580 326732 269632 326738
rect 269580 326674 269632 326680
rect 269304 326596 269356 326602
rect 269304 326538 269356 326544
rect 269488 326596 269540 326602
rect 269488 326538 269540 326544
rect 268568 326392 268620 326398
rect 268568 326334 268620 326340
rect 269212 326324 269264 326330
rect 269212 326266 269264 326272
rect 268384 280832 268436 280838
rect 268384 280774 268436 280780
rect 269224 228410 269252 326266
rect 269316 229770 269344 326538
rect 269592 326482 269620 326674
rect 269408 326454 269620 326482
rect 269408 260166 269436 326454
rect 269488 326392 269540 326398
rect 269488 326334 269540 326340
rect 269396 260160 269448 260166
rect 269396 260102 269448 260108
rect 269304 229764 269356 229770
rect 269304 229706 269356 229712
rect 269212 228404 269264 228410
rect 269212 228346 269264 228352
rect 269500 36582 269528 326334
rect 269684 326262 269712 338014
rect 269764 336048 269816 336054
rect 269764 335990 269816 335996
rect 269672 326256 269724 326262
rect 269672 326198 269724 326204
rect 269776 287706 269804 335990
rect 269960 326398 269988 338014
rect 269948 326392 270000 326398
rect 269948 326334 270000 326340
rect 270236 326330 270264 338014
rect 270224 326324 270276 326330
rect 270224 326266 270276 326272
rect 270512 313954 270540 338014
rect 270788 331214 270816 338014
rect 271064 336054 271092 338014
rect 271144 336728 271196 336734
rect 271144 336670 271196 336676
rect 271052 336048 271104 336054
rect 271052 335990 271104 335996
rect 270604 331186 270816 331214
rect 270500 313948 270552 313954
rect 270500 313890 270552 313896
rect 269764 287700 269816 287706
rect 269764 287642 269816 287648
rect 270604 246362 270632 331186
rect 270868 326392 270920 326398
rect 270868 326334 270920 326340
rect 270776 326324 270828 326330
rect 270776 326266 270828 326272
rect 270788 316674 270816 326266
rect 270776 316668 270828 316674
rect 270776 316610 270828 316616
rect 270592 246356 270644 246362
rect 270592 246298 270644 246304
rect 270880 244934 270908 326334
rect 270868 244928 270920 244934
rect 270868 244870 270920 244876
rect 271156 39370 271184 336670
rect 271236 335844 271288 335850
rect 271236 335786 271288 335792
rect 271248 254590 271276 335786
rect 271340 326330 271368 338014
rect 271616 326398 271644 338014
rect 271604 326392 271656 326398
rect 271604 326334 271656 326340
rect 271328 326324 271380 326330
rect 271328 326266 271380 326272
rect 271984 269822 272012 338014
rect 272168 336666 272196 338014
rect 272156 336660 272208 336666
rect 272156 336602 272208 336608
rect 272444 335354 272472 338014
rect 272076 335326 272472 335354
rect 272076 315314 272104 335326
rect 272064 315308 272116 315314
rect 272064 315250 272116 315256
rect 272720 311894 272748 338014
rect 272996 335850 273024 338014
rect 273272 336734 273300 338014
rect 273260 336728 273312 336734
rect 273260 336670 273312 336676
rect 272984 335844 273036 335850
rect 272984 335786 273036 335792
rect 273444 330472 273496 330478
rect 273444 330414 273496 330420
rect 273352 330404 273404 330410
rect 273352 330346 273404 330352
rect 272168 311866 272748 311894
rect 271972 269816 272024 269822
rect 271972 269758 272024 269764
rect 271236 254584 271288 254590
rect 271236 254526 271288 254532
rect 272168 227050 272196 311866
rect 272156 227044 272208 227050
rect 272156 226986 272208 226992
rect 273364 225622 273392 330346
rect 273456 243574 273484 330414
rect 273548 268394 273576 338014
rect 273824 316034 273852 338014
rect 273904 336728 273956 336734
rect 273904 336670 273956 336676
rect 273640 316006 273852 316034
rect 273536 268388 273588 268394
rect 273536 268330 273588 268336
rect 273444 243568 273496 243574
rect 273444 243510 273496 243516
rect 273352 225616 273404 225622
rect 273352 225558 273404 225564
rect 271144 39364 271196 39370
rect 271144 39306 271196 39312
rect 269488 36576 269540 36582
rect 269488 36518 269540 36524
rect 269120 18692 269172 18698
rect 269120 18634 269172 18640
rect 269132 16574 269160 18634
rect 269132 16546 270080 16574
rect 268844 7608 268896 7614
rect 268844 7550 268896 7556
rect 268108 3392 268160 3398
rect 268108 3334 268160 3340
rect 268856 480 268884 7550
rect 270052 480 270080 16546
rect 273352 14612 273404 14618
rect 273352 14554 273404 14560
rect 270776 10464 270828 10470
rect 270776 10406 270828 10412
rect 265318 354 265430 480
rect 265176 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270788 354 270816 10406
rect 272432 4888 272484 4894
rect 272432 4830 272484 4836
rect 272444 480 272472 4830
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273364 354 273392 14554
rect 273640 10334 273668 316006
rect 273916 309806 273944 336670
rect 274100 330478 274128 338014
rect 274088 330472 274140 330478
rect 274088 330414 274140 330420
rect 274376 330410 274404 338014
rect 274824 330472 274876 330478
rect 274824 330414 274876 330420
rect 274364 330404 274416 330410
rect 274364 330346 274416 330352
rect 274732 330404 274784 330410
rect 274732 330346 274784 330352
rect 273904 309800 273956 309806
rect 273904 309742 273956 309748
rect 274744 242214 274772 330346
rect 274836 284986 274864 330414
rect 274928 307086 274956 338014
rect 275020 338014 275080 338042
rect 275204 338014 275356 338042
rect 275480 338014 275632 338042
rect 275756 338014 275908 338042
rect 276124 338014 276184 338042
rect 276308 338014 276460 338042
rect 276584 338014 276736 338042
rect 276860 338014 277012 338042
rect 277136 338014 277288 338042
rect 277504 338014 277564 338042
rect 277780 338014 277840 338042
rect 277964 338014 278116 338042
rect 278240 338014 278392 338042
rect 278516 338014 278668 338042
rect 278944 338014 279096 338042
rect 275020 336734 275048 338014
rect 275008 336728 275060 336734
rect 275008 336670 275060 336676
rect 275204 316034 275232 338014
rect 275284 335708 275336 335714
rect 275284 335650 275336 335656
rect 275020 316006 275232 316034
rect 274916 307080 274968 307086
rect 274916 307022 274968 307028
rect 274824 284980 274876 284986
rect 274824 284922 274876 284928
rect 274732 242208 274784 242214
rect 274732 242150 274784 242156
rect 275020 42090 275048 316006
rect 275296 253230 275324 335650
rect 275480 330478 275508 338014
rect 275468 330472 275520 330478
rect 275468 330414 275520 330420
rect 275756 330410 275784 338014
rect 275744 330404 275796 330410
rect 275744 330346 275796 330352
rect 276124 275330 276152 338014
rect 276308 335714 276336 338014
rect 276296 335708 276348 335714
rect 276296 335650 276348 335656
rect 276584 335354 276612 338014
rect 276216 335326 276612 335354
rect 276216 319462 276244 335326
rect 276204 319456 276256 319462
rect 276204 319398 276256 319404
rect 276860 316034 276888 338014
rect 277136 327758 277164 338014
rect 277400 330472 277452 330478
rect 277400 330414 277452 330420
rect 277124 327752 277176 327758
rect 277124 327694 277176 327700
rect 276308 316006 276888 316034
rect 276112 275324 276164 275330
rect 276112 275266 276164 275272
rect 275284 253224 275336 253230
rect 275284 253166 275336 253172
rect 276308 221474 276336 316006
rect 276296 221468 276348 221474
rect 276296 221410 276348 221416
rect 275008 42084 275060 42090
rect 275008 42026 275060 42032
rect 277412 15978 277440 330414
rect 277400 15972 277452 15978
rect 277400 15914 277452 15920
rect 277504 15910 277532 338014
rect 277676 329860 277728 329866
rect 277676 329802 277728 329808
rect 277584 329316 277636 329322
rect 277584 329258 277636 329264
rect 277596 220114 277624 329258
rect 277688 283626 277716 329802
rect 277780 304298 277808 338014
rect 277964 329866 277992 338014
rect 278240 330478 278268 338014
rect 278228 330472 278280 330478
rect 278228 330414 278280 330420
rect 277952 329860 278004 329866
rect 277952 329802 278004 329808
rect 278516 329322 278544 338014
rect 278872 336728 278924 336734
rect 278872 336670 278924 336676
rect 278504 329316 278556 329322
rect 278504 329258 278556 329264
rect 277768 304292 277820 304298
rect 277768 304234 277820 304240
rect 277676 283620 277728 283626
rect 277676 283562 277728 283568
rect 278884 239426 278912 336670
rect 278964 330540 279016 330546
rect 278964 330482 279016 330488
rect 278976 286346 279004 330482
rect 279068 318102 279096 338014
rect 279160 338014 279220 338042
rect 279344 338014 279496 338042
rect 279620 338014 279772 338042
rect 279896 338014 280048 338042
rect 280264 338014 280324 338042
rect 280448 338014 280600 338042
rect 280724 338014 280876 338042
rect 281000 338014 281152 338042
rect 281276 338014 281428 338042
rect 279160 336734 279188 338014
rect 279148 336728 279200 336734
rect 279148 336670 279200 336676
rect 279056 318096 279108 318102
rect 279056 318038 279108 318044
rect 279344 316034 279372 338014
rect 279424 336728 279476 336734
rect 279424 336670 279476 336676
rect 279160 316006 279372 316034
rect 278964 286340 279016 286346
rect 278964 286282 279016 286288
rect 278872 239420 278924 239426
rect 278872 239362 278924 239368
rect 277584 220108 277636 220114
rect 277584 220050 277636 220056
rect 279160 47598 279188 316006
rect 279436 251870 279464 336670
rect 279620 330546 279648 338014
rect 279896 331906 279924 338014
rect 279884 331900 279936 331906
rect 279884 331842 279936 331848
rect 279608 330540 279660 330546
rect 279608 330482 279660 330488
rect 280264 273970 280292 338014
rect 280448 336734 280476 338014
rect 280436 336728 280488 336734
rect 280436 336670 280488 336676
rect 280724 335354 280752 338014
rect 280356 335326 280752 335354
rect 280356 297430 280384 335326
rect 281000 316034 281028 338014
rect 281276 330478 281304 338014
rect 281690 337770 281718 338028
rect 281828 338014 281980 338042
rect 282104 338014 282256 338042
rect 282380 338014 282532 338042
rect 282656 338014 282808 338042
rect 283084 338014 283236 338042
rect 281690 337742 281764 337770
rect 281632 330540 281684 330546
rect 281632 330482 281684 330488
rect 281264 330472 281316 330478
rect 281264 330414 281316 330420
rect 280448 316006 281028 316034
rect 280344 297424 280396 297430
rect 280344 297366 280396 297372
rect 280252 273964 280304 273970
rect 280252 273906 280304 273912
rect 279424 251864 279476 251870
rect 279424 251806 279476 251812
rect 280448 218754 280476 316006
rect 280436 218748 280488 218754
rect 280436 218690 280488 218696
rect 279148 47592 279200 47598
rect 279148 47534 279200 47540
rect 281644 16114 281672 330482
rect 281632 16108 281684 16114
rect 281632 16050 281684 16056
rect 281736 16046 281764 337742
rect 281828 272542 281856 338014
rect 282104 316034 282132 338014
rect 282182 336016 282238 336025
rect 282182 335951 282238 335960
rect 281920 316006 282132 316034
rect 281816 272536 281868 272542
rect 281816 272478 281868 272484
rect 281724 16040 281776 16046
rect 281724 15982 281776 15988
rect 277492 15904 277544 15910
rect 277492 15846 277544 15852
rect 279056 15904 279108 15910
rect 279056 15846 279108 15852
rect 278320 13252 278372 13258
rect 278320 13194 278372 13200
rect 274824 11824 274876 11830
rect 274824 11766 274876 11772
rect 273628 10328 273680 10334
rect 273628 10270 273680 10276
rect 274836 480 274864 11766
rect 276020 10328 276072 10334
rect 276020 10270 276072 10276
rect 276032 480 276060 10270
rect 277124 7676 277176 7682
rect 277124 7618 277176 7624
rect 277136 480 277164 7618
rect 278332 480 278360 13194
rect 273598 354 273710 480
rect 273364 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 354 279096 15846
rect 281920 14482 281948 316006
rect 282196 313274 282224 335951
rect 282380 330546 282408 338014
rect 282656 336122 282684 338014
rect 282644 336116 282696 336122
rect 282644 336058 282696 336064
rect 283208 335306 283236 338014
rect 283300 338014 283360 338042
rect 283484 338014 283636 338042
rect 283760 338014 283912 338042
rect 284036 338014 284188 338042
rect 284312 338014 284464 338042
rect 284588 338014 284740 338042
rect 284864 338014 285016 338042
rect 285140 338014 285292 338042
rect 285416 338014 285568 338042
rect 285784 338014 285844 338042
rect 286060 338014 286120 338042
rect 286244 338014 286396 338042
rect 286520 338014 286672 338042
rect 286796 338014 286948 338042
rect 287072 338014 287224 338042
rect 287348 338014 287500 338042
rect 287624 338014 287776 338042
rect 287900 338014 288052 338042
rect 288176 338014 288328 338042
rect 288544 338014 288604 338042
rect 288728 338014 288880 338042
rect 289004 338014 289156 338042
rect 289280 338014 289432 338042
rect 289556 338014 289708 338042
rect 289832 338014 289984 338042
rect 290108 338014 290260 338042
rect 290384 338014 290536 338042
rect 290660 338014 290812 338042
rect 290936 338014 291088 338042
rect 283196 335300 283248 335306
rect 283196 335242 283248 335248
rect 282368 330540 282420 330546
rect 282368 330482 282420 330488
rect 282920 330540 282972 330546
rect 283300 330528 283328 338014
rect 283380 335300 283432 335306
rect 283380 335242 283432 335248
rect 282920 330482 282972 330488
rect 283116 330500 283328 330528
rect 282184 313268 282236 313274
rect 282184 313210 282236 313216
rect 282932 49026 282960 330482
rect 283012 330472 283064 330478
rect 283012 330414 283064 330420
rect 283024 236706 283052 330414
rect 283116 238066 283144 330500
rect 283196 330404 283248 330410
rect 283196 330346 283248 330352
rect 283208 290494 283236 330346
rect 283392 316034 283420 335242
rect 283484 330546 283512 338014
rect 283472 330540 283524 330546
rect 283472 330482 283524 330488
rect 283760 330410 283788 338014
rect 284036 330478 284064 338014
rect 284312 336190 284340 338014
rect 284484 336728 284536 336734
rect 284484 336670 284536 336676
rect 284300 336184 284352 336190
rect 284300 336126 284352 336132
rect 284300 335980 284352 335986
rect 284300 335922 284352 335928
rect 284312 333334 284340 335922
rect 284300 333328 284352 333334
rect 284300 333270 284352 333276
rect 284392 330540 284444 330546
rect 284392 330482 284444 330488
rect 284024 330472 284076 330478
rect 284024 330414 284076 330420
rect 283748 330404 283800 330410
rect 283748 330346 283800 330352
rect 283300 316006 283420 316034
rect 283300 300150 283328 316006
rect 283288 300144 283340 300150
rect 283288 300086 283340 300092
rect 283196 290488 283248 290494
rect 283196 290430 283248 290436
rect 283104 238060 283156 238066
rect 283104 238002 283156 238008
rect 283012 236700 283064 236706
rect 283012 236642 283064 236648
rect 282920 49020 282972 49026
rect 282920 48962 282972 48968
rect 282000 15972 282052 15978
rect 282000 15914 282052 15920
rect 281908 14476 281960 14482
rect 281908 14418 281960 14424
rect 280712 10396 280764 10402
rect 280712 10338 280764 10344
rect 280724 480 280752 10338
rect 282012 6914 282040 15914
rect 284404 14550 284432 330482
rect 284496 17270 284524 336670
rect 284588 250510 284616 338014
rect 284864 336734 284892 338014
rect 284852 336728 284904 336734
rect 284852 336670 284904 336676
rect 285140 316034 285168 338014
rect 285416 330546 285444 338014
rect 285680 336048 285732 336054
rect 285680 335990 285732 335996
rect 285692 334694 285720 335990
rect 285680 334688 285732 334694
rect 285680 334630 285732 334636
rect 285404 330540 285456 330546
rect 285404 330482 285456 330488
rect 284680 316006 285168 316034
rect 284576 250504 284628 250510
rect 284576 250446 284628 250452
rect 284484 17264 284536 17270
rect 284484 17206 284536 17212
rect 284392 14544 284444 14550
rect 284392 14486 284444 14492
rect 284576 14476 284628 14482
rect 284576 14418 284628 14424
rect 283104 13184 283156 13190
rect 283104 13126 283156 13132
rect 281920 6886 282040 6914
rect 281920 480 281948 6886
rect 283116 480 283144 13126
rect 284300 3460 284352 3466
rect 284300 3402 284352 3408
rect 284312 480 284340 3402
rect 284588 490 284616 14418
rect 284680 3330 284708 316006
rect 285784 43450 285812 338014
rect 285956 330540 286008 330546
rect 285956 330482 286008 330488
rect 285864 330472 285916 330478
rect 285864 330414 285916 330420
rect 285876 51746 285904 330414
rect 285968 297498 285996 330482
rect 285956 297492 286008 297498
rect 285956 297434 286008 297440
rect 285864 51740 285916 51746
rect 285864 51682 285916 51688
rect 285956 51740 286008 51746
rect 285956 51682 286008 51688
rect 285772 43444 285824 43450
rect 285772 43386 285824 43392
rect 285680 3596 285732 3602
rect 285680 3538 285732 3544
rect 284668 3324 284720 3330
rect 284668 3266 284720 3272
rect 285692 3262 285720 3538
rect 285968 3482 285996 51682
rect 286060 3602 286088 338014
rect 286244 335986 286272 338014
rect 286232 335980 286284 335986
rect 286232 335922 286284 335928
rect 286324 335368 286376 335374
rect 286324 335310 286376 335316
rect 286336 320890 286364 335310
rect 286520 330546 286548 338014
rect 286508 330540 286560 330546
rect 286508 330482 286560 330488
rect 286796 330478 286824 338014
rect 286784 330472 286836 330478
rect 286784 330414 286836 330420
rect 287072 320890 287100 338014
rect 287348 330834 287376 338014
rect 287624 335374 287652 338014
rect 287704 336728 287756 336734
rect 287704 336670 287756 336676
rect 287612 335368 287664 335374
rect 287612 335310 287664 335316
rect 287164 330806 287376 330834
rect 286324 320884 286376 320890
rect 286324 320826 286376 320832
rect 287060 320884 287112 320890
rect 287060 320826 287112 320832
rect 287164 287774 287192 330806
rect 287336 330540 287388 330546
rect 287336 330482 287388 330488
rect 287244 320884 287296 320890
rect 287244 320826 287296 320832
rect 287256 315382 287284 320826
rect 287244 315376 287296 315382
rect 287244 315318 287296 315324
rect 287152 287768 287204 287774
rect 287152 287710 287204 287716
rect 287348 282198 287376 330482
rect 287336 282192 287388 282198
rect 287336 282134 287388 282140
rect 287716 13122 287744 336670
rect 287900 336394 287928 338014
rect 287888 336388 287940 336394
rect 287888 336330 287940 336336
rect 287796 335708 287848 335714
rect 287796 335650 287848 335656
rect 287808 312662 287836 335650
rect 288176 330546 288204 338014
rect 288164 330540 288216 330546
rect 288164 330482 288216 330488
rect 287796 312656 287848 312662
rect 287796 312598 287848 312604
rect 288544 261526 288572 338014
rect 288728 335714 288756 338014
rect 289004 336734 289032 338014
rect 288992 336728 289044 336734
rect 288992 336670 289044 336676
rect 289176 336728 289228 336734
rect 289176 336670 289228 336676
rect 288716 335708 288768 335714
rect 288716 335650 288768 335656
rect 289084 335572 289136 335578
rect 289084 335514 289136 335520
rect 288716 330540 288768 330546
rect 288716 330482 288768 330488
rect 288624 330472 288676 330478
rect 288624 330414 288676 330420
rect 288636 305726 288664 330414
rect 288624 305720 288676 305726
rect 288624 305662 288676 305668
rect 288532 261520 288584 261526
rect 288532 261462 288584 261468
rect 288728 258738 288756 330482
rect 288716 258732 288768 258738
rect 288716 258674 288768 258680
rect 289096 37942 289124 335514
rect 289188 304366 289216 336670
rect 289280 330546 289308 338014
rect 289268 330540 289320 330546
rect 289268 330482 289320 330488
rect 289556 330478 289584 338014
rect 289832 335578 289860 338014
rect 289820 335572 289872 335578
rect 289820 335514 289872 335520
rect 290108 335354 290136 338014
rect 290384 336734 290412 338014
rect 290372 336728 290424 336734
rect 290372 336670 290424 336676
rect 290016 335326 290136 335354
rect 289544 330472 289596 330478
rect 289544 330414 289596 330420
rect 289912 326188 289964 326194
rect 289912 326130 289964 326136
rect 289924 308514 289952 326130
rect 290016 322318 290044 335326
rect 290660 326194 290688 338014
rect 290648 326188 290700 326194
rect 290648 326130 290700 326136
rect 290004 322312 290056 322318
rect 290004 322254 290056 322260
rect 290936 316034 290964 338014
rect 291350 337770 291378 338028
rect 291488 338014 291640 338042
rect 291764 338014 291916 338042
rect 292040 338014 292192 338042
rect 292316 338014 292468 338042
rect 291350 337742 291424 337770
rect 291292 327072 291344 327078
rect 291292 327014 291344 327020
rect 290108 316006 290964 316034
rect 289912 308508 289964 308514
rect 289912 308450 289964 308456
rect 289176 304360 289228 304366
rect 289176 304302 289228 304308
rect 290108 257378 290136 316006
rect 291304 301578 291332 327014
rect 291396 303006 291424 337742
rect 291488 309874 291516 338014
rect 291568 330540 291620 330546
rect 291568 330482 291620 330488
rect 291476 309868 291528 309874
rect 291476 309810 291528 309816
rect 291384 303000 291436 303006
rect 291384 302942 291436 302948
rect 291292 301572 291344 301578
rect 291292 301514 291344 301520
rect 291580 276690 291608 330482
rect 291764 329118 291792 338014
rect 291844 335708 291896 335714
rect 291844 335650 291896 335656
rect 291752 329112 291804 329118
rect 291752 329054 291804 329060
rect 291568 276684 291620 276690
rect 291568 276626 291620 276632
rect 290096 257372 290148 257378
rect 290096 257314 290148 257320
rect 289084 37936 289136 37942
rect 289084 37878 289136 37884
rect 291856 22778 291884 335650
rect 292040 327078 292068 338014
rect 292316 330546 292344 338014
rect 292730 337770 292758 338028
rect 292868 338014 293020 338042
rect 293144 338014 293296 338042
rect 293420 338014 293572 338042
rect 293696 338014 293848 338042
rect 293972 338014 294124 338042
rect 294248 338014 294400 338042
rect 294524 338014 294676 338042
rect 294800 338014 294952 338042
rect 295076 338014 295228 338042
rect 295352 338014 295504 338042
rect 295628 338014 295780 338042
rect 295904 338014 296056 338042
rect 296180 338014 296332 338042
rect 296456 338014 296608 338042
rect 292730 337742 292804 337770
rect 292776 330750 292804 337742
rect 292764 330744 292816 330750
rect 292764 330686 292816 330692
rect 292868 330562 292896 338014
rect 293144 335714 293172 338014
rect 293224 336728 293276 336734
rect 293224 336670 293276 336676
rect 293132 335708 293184 335714
rect 293132 335650 293184 335656
rect 292948 330744 293000 330750
rect 292948 330686 293000 330692
rect 292304 330540 292356 330546
rect 292304 330482 292356 330488
rect 292672 330540 292724 330546
rect 292672 330482 292724 330488
rect 292776 330534 292896 330562
rect 292028 327072 292080 327078
rect 292028 327014 292080 327020
rect 292684 298858 292712 330482
rect 292776 300218 292804 330534
rect 292856 330472 292908 330478
rect 292856 330414 292908 330420
rect 292868 323678 292896 330414
rect 292856 323672 292908 323678
rect 292856 323614 292908 323620
rect 292764 300212 292816 300218
rect 292764 300154 292816 300160
rect 292672 298852 292724 298858
rect 292672 298794 292724 298800
rect 292960 256018 292988 330686
rect 292948 256012 293000 256018
rect 292948 255954 293000 255960
rect 293236 35222 293264 336670
rect 293316 335980 293368 335986
rect 293316 335922 293368 335928
rect 293328 222902 293356 335922
rect 293420 330478 293448 338014
rect 293696 330546 293724 338014
rect 293972 335986 294000 338014
rect 294248 336734 294276 338014
rect 294236 336728 294288 336734
rect 294236 336670 294288 336676
rect 294524 336054 294552 338014
rect 294512 336048 294564 336054
rect 294512 335990 294564 335996
rect 293960 335980 294012 335986
rect 293960 335922 294012 335928
rect 293684 330540 293736 330546
rect 293684 330482 293736 330488
rect 293408 330472 293460 330478
rect 293408 330414 293460 330420
rect 294800 327826 294828 338014
rect 294788 327820 294840 327826
rect 294788 327762 294840 327768
rect 295076 316034 295104 338014
rect 295352 325038 295380 338014
rect 295628 330426 295656 338014
rect 295444 330398 295656 330426
rect 295340 325032 295392 325038
rect 295340 324974 295392 324980
rect 294156 316006 295104 316034
rect 294156 275398 294184 316006
rect 295444 296070 295472 330398
rect 295904 316034 295932 338014
rect 296180 336462 296208 338014
rect 296168 336456 296220 336462
rect 296168 336398 296220 336404
rect 296456 336326 296484 338014
rect 296870 337770 296898 338028
rect 297008 338014 297160 338042
rect 297284 338014 297436 338042
rect 297560 338014 297712 338042
rect 297836 338014 297988 338042
rect 298112 338014 298264 338042
rect 298388 338014 298540 338042
rect 298664 338014 298816 338042
rect 298940 338014 299092 338042
rect 299216 338014 299368 338042
rect 299492 338014 299644 338042
rect 299860 338014 299920 338042
rect 300044 338014 300196 338042
rect 300320 338014 300472 338042
rect 300596 338014 300748 338042
rect 300964 338014 301024 338042
rect 301148 338014 301300 338042
rect 301424 338014 301576 338042
rect 301700 338014 301852 338042
rect 301976 338014 302128 338042
rect 296870 337742 296944 337770
rect 296812 336728 296864 336734
rect 296812 336670 296864 336676
rect 296444 336320 296496 336326
rect 296444 336262 296496 336268
rect 295984 336116 296036 336122
rect 295984 336058 296036 336064
rect 295628 316006 295932 316034
rect 295432 296064 295484 296070
rect 295432 296006 295484 296012
rect 294144 275392 294196 275398
rect 294144 275334 294196 275340
rect 295628 274038 295656 316006
rect 295616 274032 295668 274038
rect 295616 273974 295668 273980
rect 293316 222896 293368 222902
rect 293316 222838 293368 222844
rect 293224 35216 293276 35222
rect 293224 35158 293276 35164
rect 291844 22772 291896 22778
rect 291844 22714 291896 22720
rect 292580 22772 292632 22778
rect 292580 22714 292632 22720
rect 292592 16574 292620 22714
rect 295340 17264 295392 17270
rect 295340 17206 295392 17212
rect 295352 16574 295380 17206
rect 292592 16546 293264 16574
rect 295352 16546 295656 16574
rect 287704 13116 287756 13122
rect 287704 13058 287756 13064
rect 292580 7812 292632 7818
rect 292580 7754 292632 7760
rect 288992 6316 289044 6322
rect 288992 6258 289044 6264
rect 286048 3596 286100 3602
rect 286048 3538 286100 3544
rect 285968 3454 286640 3482
rect 285680 3256 285732 3262
rect 285680 3198 285732 3204
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 284588 462 284984 490
rect 286612 480 286640 3454
rect 287796 3324 287848 3330
rect 287796 3266 287848 3272
rect 287808 480 287836 3266
rect 289004 480 289032 6258
rect 290188 4956 290240 4962
rect 290188 4898 290240 4904
rect 290200 480 290228 4898
rect 291384 3596 291436 3602
rect 291384 3538 291436 3544
rect 291396 480 291424 3538
rect 292592 480 292620 7754
rect 284956 354 284984 462
rect 285374 354 285486 480
rect 284956 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 294880 3664 294932 3670
rect 294880 3606 294932 3612
rect 294892 480 294920 3606
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 295628 354 295656 16546
rect 295996 5030 296024 336058
rect 296168 335504 296220 335510
rect 296168 335446 296220 335452
rect 296076 335436 296128 335442
rect 296076 335378 296128 335384
rect 296088 18630 296116 335378
rect 296180 24138 296208 335446
rect 296260 335368 296312 335374
rect 296260 335310 296312 335316
rect 296272 323746 296300 335310
rect 296260 323740 296312 323746
rect 296260 323682 296312 323688
rect 296720 294636 296772 294642
rect 296720 294578 296772 294584
rect 296168 24132 296220 24138
rect 296168 24074 296220 24080
rect 296076 18624 296128 18630
rect 296076 18566 296128 18572
rect 296732 16574 296760 294578
rect 296824 271182 296852 336670
rect 296916 272610 296944 337742
rect 297008 335374 297036 338014
rect 297180 336048 297232 336054
rect 297180 335990 297232 335996
rect 296996 335368 297048 335374
rect 296996 335310 297048 335316
rect 296996 330540 297048 330546
rect 296996 330482 297048 330488
rect 297008 322386 297036 330482
rect 297192 325694 297220 335990
rect 297284 335442 297312 338014
rect 297560 336734 297588 338014
rect 297548 336728 297600 336734
rect 297548 336670 297600 336676
rect 297548 336184 297600 336190
rect 297548 336126 297600 336132
rect 297456 335640 297508 335646
rect 297456 335582 297508 335588
rect 297272 335436 297324 335442
rect 297272 335378 297324 335384
rect 297192 325666 297404 325694
rect 296996 322380 297048 322386
rect 296996 322322 297048 322328
rect 296904 272604 296956 272610
rect 296904 272546 296956 272552
rect 296812 271176 296864 271182
rect 296812 271118 296864 271124
rect 296732 16546 297312 16574
rect 295984 5024 296036 5030
rect 295984 4966 296036 4972
rect 297284 480 297312 16546
rect 297376 6322 297404 325666
rect 297468 294710 297496 335582
rect 297560 320958 297588 336126
rect 297836 330546 297864 338014
rect 298112 335646 298140 338014
rect 298100 335640 298152 335646
rect 298100 335582 298152 335588
rect 298388 335510 298416 338014
rect 298664 336190 298692 338014
rect 298744 336728 298796 336734
rect 298744 336670 298796 336676
rect 298652 336184 298704 336190
rect 298652 336126 298704 336132
rect 298376 335504 298428 335510
rect 298376 335446 298428 335452
rect 297824 330540 297876 330546
rect 297824 330482 297876 330488
rect 298192 330540 298244 330546
rect 298192 330482 298244 330488
rect 297548 320952 297600 320958
rect 297548 320894 297600 320900
rect 298204 307154 298232 330482
rect 298284 330472 298336 330478
rect 298284 330414 298336 330420
rect 298192 307148 298244 307154
rect 298192 307090 298244 307096
rect 297456 294704 297508 294710
rect 297456 294646 297508 294652
rect 298296 269890 298324 330414
rect 298284 269884 298336 269890
rect 298284 269826 298336 269832
rect 298756 268462 298784 336670
rect 298940 330546 298968 338014
rect 298928 330540 298980 330546
rect 298928 330482 298980 330488
rect 299216 330478 299244 338014
rect 299204 330472 299256 330478
rect 299204 330414 299256 330420
rect 299492 326466 299520 338014
rect 299860 330562 299888 338014
rect 300044 336734 300072 338014
rect 300032 336728 300084 336734
rect 300032 336670 300084 336676
rect 300124 336184 300176 336190
rect 300124 336126 300176 336132
rect 299584 330534 299888 330562
rect 299480 326460 299532 326466
rect 299480 326402 299532 326408
rect 299584 291922 299612 330534
rect 299848 330404 299900 330410
rect 299848 330346 299900 330352
rect 299664 330336 299716 330342
rect 299664 330278 299716 330284
rect 299676 318170 299704 330278
rect 299664 318164 299716 318170
rect 299664 318106 299716 318112
rect 299664 292052 299716 292058
rect 299664 291994 299716 292000
rect 299572 291916 299624 291922
rect 299572 291858 299624 291864
rect 298744 268456 298796 268462
rect 298744 268398 298796 268404
rect 299480 18624 299532 18630
rect 299480 18566 299532 18572
rect 299492 6914 299520 18566
rect 299676 16574 299704 291994
rect 299860 25566 299888 330346
rect 299848 25560 299900 25566
rect 299848 25502 299900 25508
rect 299676 16546 299796 16574
rect 299768 6914 299796 16546
rect 300136 13258 300164 336126
rect 300320 330342 300348 338014
rect 300596 330410 300624 338014
rect 300860 336728 300912 336734
rect 300860 336670 300912 336676
rect 300584 330404 300636 330410
rect 300584 330346 300636 330352
rect 300308 330336 300360 330342
rect 300308 330278 300360 330284
rect 300872 327894 300900 336670
rect 300860 327888 300912 327894
rect 300860 327830 300912 327836
rect 300964 265674 300992 338014
rect 301148 336734 301176 338014
rect 301424 336818 301452 338014
rect 301240 336790 301452 336818
rect 301136 336728 301188 336734
rect 301136 336670 301188 336676
rect 301240 335354 301268 336790
rect 301700 336682 301728 338014
rect 301056 335326 301268 335354
rect 301424 336654 301728 336682
rect 301056 290562 301084 335326
rect 301136 330540 301188 330546
rect 301136 330482 301188 330488
rect 301148 316810 301176 330482
rect 301136 316804 301188 316810
rect 301136 316746 301188 316752
rect 301424 316034 301452 336654
rect 301504 336456 301556 336462
rect 301504 336398 301556 336404
rect 301240 316006 301452 316034
rect 301044 290556 301096 290562
rect 301044 290498 301096 290504
rect 300952 265668 301004 265674
rect 300952 265610 301004 265616
rect 301240 264246 301268 316006
rect 301228 264240 301280 264246
rect 301228 264182 301280 264188
rect 300124 13252 300176 13258
rect 300124 13194 300176 13200
rect 301516 7750 301544 336398
rect 301976 330546 302004 338014
rect 302390 337770 302418 338028
rect 302528 338014 302680 338042
rect 302804 338014 302956 338042
rect 303080 338014 303232 338042
rect 303356 338014 303508 338042
rect 303784 338014 303936 338042
rect 302390 337742 302464 337770
rect 302240 336728 302292 336734
rect 302240 336670 302292 336676
rect 301964 330540 302016 330546
rect 301964 330482 302016 330488
rect 302252 26926 302280 336670
rect 302332 326460 302384 326466
rect 302332 326402 302384 326408
rect 302344 262954 302372 326402
rect 302436 289202 302464 337742
rect 302528 336734 302556 338014
rect 302516 336728 302568 336734
rect 302516 336670 302568 336676
rect 302804 335354 302832 338014
rect 302528 335326 302832 335354
rect 302884 335368 302936 335374
rect 302528 314022 302556 335326
rect 302884 335310 302936 335316
rect 302608 326392 302660 326398
rect 302608 326334 302660 326340
rect 302620 318238 302648 326334
rect 302608 318232 302660 318238
rect 302608 318174 302660 318180
rect 302516 314016 302568 314022
rect 302516 313958 302568 313964
rect 302424 289196 302476 289202
rect 302424 289138 302476 289144
rect 302332 262948 302384 262954
rect 302332 262890 302384 262896
rect 302896 29646 302924 335310
rect 303080 326398 303108 338014
rect 303356 326466 303384 338014
rect 303620 336728 303672 336734
rect 303620 336670 303672 336676
rect 303528 336660 303580 336666
rect 303528 336602 303580 336608
rect 303540 334830 303568 336602
rect 303528 334824 303580 334830
rect 303528 334766 303580 334772
rect 303632 326534 303660 336670
rect 303620 326528 303672 326534
rect 303620 326470 303672 326476
rect 303344 326460 303396 326466
rect 303344 326402 303396 326408
rect 303068 326392 303120 326398
rect 303068 326334 303120 326340
rect 303804 326392 303856 326398
rect 303804 326334 303856 326340
rect 303712 326324 303764 326330
rect 303712 326266 303764 326272
rect 303620 318096 303672 318102
rect 303620 318038 303672 318044
rect 302884 29640 302936 29646
rect 302884 29582 302936 29588
rect 302240 26920 302292 26926
rect 302240 26862 302292 26868
rect 303632 16574 303660 318038
rect 303724 21418 303752 326266
rect 303816 304434 303844 326334
rect 303908 319530 303936 338014
rect 304000 338014 304060 338042
rect 304184 338014 304336 338042
rect 304460 338014 304612 338042
rect 304736 338014 304888 338042
rect 305012 338014 305164 338042
rect 305380 338014 305440 338042
rect 305564 338014 305716 338042
rect 305840 338014 305992 338042
rect 306116 338014 306268 338042
rect 304000 336734 304028 338014
rect 303988 336728 304040 336734
rect 303988 336670 304040 336676
rect 303988 326460 304040 326466
rect 303988 326402 304040 326408
rect 303896 319524 303948 319530
rect 303896 319466 303948 319472
rect 304000 311234 304028 326402
rect 304184 326398 304212 338014
rect 304264 336320 304316 336326
rect 304264 336262 304316 336268
rect 304172 326392 304224 326398
rect 304172 326334 304224 326340
rect 303988 311228 304040 311234
rect 303988 311170 304040 311176
rect 303804 304428 303856 304434
rect 303804 304370 303856 304376
rect 303712 21412 303764 21418
rect 303712 21354 303764 21360
rect 303632 16546 303936 16574
rect 303160 13116 303212 13122
rect 303160 13058 303212 13064
rect 301504 7744 301556 7750
rect 301504 7686 301556 7692
rect 299492 6886 299704 6914
rect 299768 6886 300808 6914
rect 297364 6316 297416 6322
rect 297364 6258 297416 6264
rect 298468 3732 298520 3738
rect 298468 3674 298520 3680
rect 298480 480 298508 3674
rect 299676 480 299704 6886
rect 300780 480 300808 6886
rect 301964 3800 302016 3806
rect 301964 3742 302016 3748
rect 301976 480 302004 3742
rect 303172 480 303200 13058
rect 296046 354 296158 480
rect 295628 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 304276 15978 304304 336262
rect 304460 326466 304488 338014
rect 304448 326460 304500 326466
rect 304448 326402 304500 326408
rect 304736 326330 304764 338014
rect 305012 334762 305040 338014
rect 305000 334756 305052 334762
rect 305000 334698 305052 334704
rect 305380 331974 305408 338014
rect 305564 335354 305592 338014
rect 305736 336592 305788 336598
rect 305736 336534 305788 336540
rect 305644 336388 305696 336394
rect 305644 336330 305696 336336
rect 305472 335326 305592 335354
rect 305368 331968 305420 331974
rect 305368 331910 305420 331916
rect 305472 331214 305500 335326
rect 305104 331186 305500 331214
rect 304724 326324 304776 326330
rect 304724 326266 304776 326272
rect 305104 286414 305132 331186
rect 305184 326460 305236 326466
rect 305184 326402 305236 326408
rect 305196 309942 305224 326402
rect 305276 326392 305328 326398
rect 305276 326334 305328 326340
rect 305184 309936 305236 309942
rect 305184 309878 305236 309884
rect 305092 286408 305144 286414
rect 305092 286350 305144 286356
rect 305288 28286 305316 326334
rect 305276 28280 305328 28286
rect 305276 28222 305328 28228
rect 304264 15972 304316 15978
rect 304264 15914 304316 15920
rect 305656 14482 305684 336330
rect 305748 319598 305776 336534
rect 305840 326398 305868 338014
rect 306116 326466 306144 338014
rect 306530 337770 306558 338028
rect 306668 338014 306820 338042
rect 306944 338014 307096 338042
rect 307220 338014 307372 338042
rect 307496 338014 307648 338042
rect 307772 338014 307924 338042
rect 308048 338014 308200 338042
rect 308324 338014 308476 338042
rect 308600 338014 308752 338042
rect 308876 338014 309028 338042
rect 309304 338014 309456 338042
rect 306530 337742 306604 337770
rect 306104 326460 306156 326466
rect 306104 326402 306156 326408
rect 305828 326392 305880 326398
rect 305828 326334 305880 326340
rect 306472 323740 306524 323746
rect 306472 323682 306524 323688
rect 305736 319592 305788 319598
rect 305736 319534 305788 319540
rect 306484 293282 306512 323682
rect 306576 315450 306604 337742
rect 306668 335374 306696 338014
rect 306656 335368 306708 335374
rect 306656 335310 306708 335316
rect 306944 330614 306972 338014
rect 307024 336524 307076 336530
rect 307024 336466 307076 336472
rect 306932 330608 306984 330614
rect 306932 330550 306984 330556
rect 306656 326392 306708 326398
rect 306656 326334 306708 326340
rect 306564 315444 306616 315450
rect 306564 315386 306616 315392
rect 306472 293276 306524 293282
rect 306472 293218 306524 293224
rect 306668 188358 306696 326334
rect 306656 188352 306708 188358
rect 306656 188294 306708 188300
rect 305644 14476 305696 14482
rect 305644 14418 305696 14424
rect 306380 14476 306432 14482
rect 306380 14418 306432 14424
rect 305552 3868 305604 3874
rect 305552 3810 305604 3816
rect 305564 480 305592 3810
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306392 354 306420 14418
rect 307036 13190 307064 336466
rect 307220 323746 307248 338014
rect 307496 326398 307524 338014
rect 307772 336258 307800 338014
rect 307760 336252 307812 336258
rect 307760 336194 307812 336200
rect 308048 335354 308076 338014
rect 307956 335326 308076 335354
rect 307484 326392 307536 326398
rect 307484 326334 307536 326340
rect 307852 326392 307904 326398
rect 307852 326334 307904 326340
rect 307208 323740 307260 323746
rect 307208 323682 307260 323688
rect 307864 303074 307892 326334
rect 307956 316878 307984 335326
rect 308324 326398 308352 338014
rect 308600 333402 308628 338014
rect 308588 333396 308640 333402
rect 308588 333338 308640 333344
rect 308312 326392 308364 326398
rect 308312 326334 308364 326340
rect 307944 316872 307996 316878
rect 307944 316814 307996 316820
rect 308876 316034 308904 338014
rect 309324 326460 309376 326466
rect 309324 326402 309376 326408
rect 309232 325372 309284 325378
rect 309232 325314 309284 325320
rect 308048 316006 308904 316034
rect 307852 303068 307904 303074
rect 307852 303010 307904 303016
rect 307760 285184 307812 285190
rect 307760 285126 307812 285132
rect 307772 16574 307800 285126
rect 308048 285054 308076 316006
rect 308036 285048 308088 285054
rect 308036 284990 308088 284996
rect 309244 283694 309272 325314
rect 309336 308582 309364 326402
rect 309428 312730 309456 338014
rect 309566 337770 309594 338028
rect 309704 338014 309856 338042
rect 309980 338014 310132 338042
rect 310256 338014 310408 338042
rect 310624 338014 310684 338042
rect 310900 338014 310960 338042
rect 311084 338014 311236 338042
rect 311360 338014 311512 338042
rect 311636 338014 311788 338042
rect 311912 338014 312064 338042
rect 312188 338014 312340 338042
rect 312464 338014 312616 338042
rect 312740 338014 312892 338042
rect 313016 338014 313168 338042
rect 313384 338014 313444 338042
rect 313568 338014 313720 338042
rect 313844 338014 313996 338042
rect 314120 338014 314272 338042
rect 314396 338014 314548 338042
rect 309566 337742 309640 337770
rect 309612 329186 309640 337742
rect 309600 329180 309652 329186
rect 309600 329122 309652 329128
rect 309508 326392 309560 326398
rect 309508 326334 309560 326340
rect 309416 312724 309468 312730
rect 309416 312666 309468 312672
rect 309324 308576 309376 308582
rect 309324 308518 309376 308524
rect 309232 283688 309284 283694
rect 309232 283630 309284 283636
rect 309520 31074 309548 326334
rect 309704 325378 309732 338014
rect 309876 336728 309928 336734
rect 309876 336670 309928 336676
rect 309784 336252 309836 336258
rect 309784 336194 309836 336200
rect 309692 325372 309744 325378
rect 309692 325314 309744 325320
rect 309508 31068 309560 31074
rect 309508 31010 309560 31016
rect 307772 16546 307984 16574
rect 307024 13184 307076 13190
rect 307024 13126 307076 13132
rect 307956 480 307984 16546
rect 309796 10470 309824 336194
rect 309888 323814 309916 336670
rect 309980 326398 310008 338014
rect 310256 326466 310284 338014
rect 310244 326460 310296 326466
rect 310244 326402 310296 326408
rect 309968 326392 310020 326398
rect 309968 326334 310020 326340
rect 310624 326262 310652 338014
rect 310900 326346 310928 338014
rect 310716 326318 310928 326346
rect 310612 326256 310664 326262
rect 310612 326198 310664 326204
rect 310612 324284 310664 324290
rect 310612 324226 310664 324232
rect 309876 323808 309928 323814
rect 309876 323750 309928 323756
rect 310624 280906 310652 324226
rect 310716 301646 310744 326318
rect 310796 326256 310848 326262
rect 310796 326198 310848 326204
rect 310888 326256 310940 326262
rect 310888 326198 310940 326204
rect 310808 314090 310836 326198
rect 310796 314084 310848 314090
rect 310796 314026 310848 314032
rect 310704 301640 310756 301646
rect 310704 301582 310756 301588
rect 310612 280900 310664 280906
rect 310612 280842 310664 280848
rect 310900 267034 310928 326198
rect 311084 325106 311112 338014
rect 311164 335504 311216 335510
rect 311164 335446 311216 335452
rect 311072 325100 311124 325106
rect 311072 325042 311124 325048
rect 310888 267028 310940 267034
rect 310888 266970 310940 266976
rect 310520 21412 310572 21418
rect 310520 21354 310572 21360
rect 309876 10532 309928 10538
rect 309876 10474 309928 10480
rect 309784 10464 309836 10470
rect 309784 10406 309836 10412
rect 309888 6914 309916 10474
rect 309796 6886 309916 6914
rect 310532 6914 310560 21354
rect 311176 9110 311204 335446
rect 311360 324290 311388 338014
rect 311636 326262 311664 338014
rect 311912 336666 311940 338014
rect 311900 336660 311952 336666
rect 311900 336602 311952 336608
rect 312188 335354 312216 338014
rect 312096 335326 312216 335354
rect 311992 328364 312044 328370
rect 311992 328306 312044 328312
rect 311624 326256 311676 326262
rect 311624 326198 311676 326204
rect 311348 324284 311400 324290
rect 311348 324226 311400 324232
rect 312004 279546 312032 328306
rect 312096 311302 312124 335326
rect 312464 316034 312492 338014
rect 312740 336734 312768 338014
rect 312728 336728 312780 336734
rect 312728 336670 312780 336676
rect 313016 328370 313044 338014
rect 313004 328364 313056 328370
rect 313004 328306 313056 328312
rect 312188 316006 312492 316034
rect 312084 311296 312136 311302
rect 312084 311238 312136 311244
rect 311992 279540 312044 279546
rect 311992 279482 312044 279488
rect 312188 240786 312216 316006
rect 313384 260234 313412 338014
rect 313464 330472 313516 330478
rect 313464 330414 313516 330420
rect 313476 307222 313504 330414
rect 313568 322454 313596 338014
rect 313844 332042 313872 338014
rect 313924 335368 313976 335374
rect 313924 335310 313976 335316
rect 313832 332036 313884 332042
rect 313832 331978 313884 331984
rect 313648 330540 313700 330546
rect 313648 330482 313700 330488
rect 313556 322448 313608 322454
rect 313556 322390 313608 322396
rect 313464 307216 313516 307222
rect 313464 307158 313516 307164
rect 313372 260228 313424 260234
rect 313372 260170 313424 260176
rect 312176 240780 312228 240786
rect 312176 240722 312228 240728
rect 313660 33794 313688 330482
rect 313648 33788 313700 33794
rect 313648 33730 313700 33736
rect 311164 9104 311216 9110
rect 311164 9046 311216 9052
rect 310532 6886 311480 6914
rect 309048 3936 309100 3942
rect 309048 3878 309100 3884
rect 309060 480 309088 3878
rect 306718 354 306830 480
rect 306392 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 6886
rect 311452 480 311480 6886
rect 313832 5024 313884 5030
rect 313832 4966 313884 4972
rect 312636 4004 312688 4010
rect 312636 3946 312688 3952
rect 312648 480 312676 3946
rect 313844 480 313872 4966
rect 313936 4826 313964 335310
rect 314120 330546 314148 338014
rect 314108 330540 314160 330546
rect 314108 330482 314160 330488
rect 314396 330478 314424 338014
rect 314810 337770 314838 338028
rect 314948 338014 315100 338042
rect 315224 338014 315376 338042
rect 315500 338014 315652 338042
rect 315776 338014 315928 338042
rect 316052 338014 316204 338042
rect 316328 338014 316480 338042
rect 316604 338014 316756 338042
rect 316880 338014 317032 338042
rect 317156 338014 317308 338042
rect 314810 337742 314884 337770
rect 314384 330472 314436 330478
rect 314384 330414 314436 330420
rect 314752 327752 314804 327758
rect 314752 327694 314804 327700
rect 314660 278248 314712 278254
rect 314660 278190 314712 278196
rect 313924 4820 313976 4826
rect 313924 4762 313976 4768
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314672 354 314700 278190
rect 314764 166326 314792 327694
rect 314856 305794 314884 337742
rect 314948 333470 314976 338014
rect 315224 335354 315252 338014
rect 315304 335708 315356 335714
rect 315304 335650 315356 335656
rect 315040 335326 315252 335354
rect 314936 333464 314988 333470
rect 314936 333406 314988 333412
rect 315040 330562 315068 335326
rect 314948 330534 315068 330562
rect 314948 321026 314976 330534
rect 315028 330472 315080 330478
rect 315028 330414 315080 330420
rect 314936 321020 314988 321026
rect 314936 320962 314988 320968
rect 314844 305788 314896 305794
rect 314844 305730 314896 305736
rect 315040 278118 315068 330414
rect 315028 278112 315080 278118
rect 315028 278054 315080 278060
rect 314752 166320 314804 166326
rect 314752 166262 314804 166268
rect 315316 6186 315344 335650
rect 315500 330478 315528 338014
rect 315488 330472 315540 330478
rect 315488 330414 315540 330420
rect 315776 327758 315804 338014
rect 316052 336598 316080 338014
rect 316040 336592 316092 336598
rect 316040 336534 316092 336540
rect 316328 330682 316356 338014
rect 316316 330676 316368 330682
rect 316316 330618 316368 330624
rect 315764 327752 315816 327758
rect 315764 327694 315816 327700
rect 316604 316034 316632 338014
rect 316684 336592 316736 336598
rect 316684 336534 316736 336540
rect 316236 316006 316632 316034
rect 316236 297566 316264 316006
rect 316224 297560 316276 297566
rect 316224 297502 316276 297508
rect 316696 15910 316724 336534
rect 316880 335374 316908 338014
rect 317156 335714 317184 338014
rect 317570 337770 317598 338028
rect 317708 338014 317860 338042
rect 317984 338014 318136 338042
rect 318260 338014 318412 338042
rect 318536 338014 318688 338042
rect 317570 337742 317644 337770
rect 317144 335708 317196 335714
rect 317144 335650 317196 335656
rect 316868 335368 316920 335374
rect 316868 335310 316920 335316
rect 317512 330472 317564 330478
rect 317512 330414 317564 330420
rect 316684 15904 316736 15910
rect 316684 15846 316736 15852
rect 317524 8974 317552 330414
rect 317616 17338 317644 337742
rect 317708 336462 317736 338014
rect 317696 336456 317748 336462
rect 317696 336398 317748 336404
rect 317984 335510 318012 338014
rect 318064 336660 318116 336666
rect 318064 336602 318116 336608
rect 317972 335504 318024 335510
rect 317972 335446 318024 335452
rect 317696 330540 317748 330546
rect 317696 330482 317748 330488
rect 317604 17332 317656 17338
rect 317604 17274 317656 17280
rect 317512 8968 317564 8974
rect 317512 8910 317564 8916
rect 317708 6254 317736 330482
rect 317696 6248 317748 6254
rect 317696 6190 317748 6196
rect 315304 6180 315356 6186
rect 315304 6122 315356 6128
rect 318076 4894 318104 336602
rect 318260 330546 318288 338014
rect 318248 330540 318300 330546
rect 318248 330482 318300 330488
rect 318536 330478 318564 338014
rect 318950 337770 318978 338028
rect 319088 338014 319240 338042
rect 319364 338014 319516 338042
rect 319640 338014 319792 338042
rect 319916 338014 320068 338042
rect 320192 338014 320344 338042
rect 320468 338014 320620 338042
rect 320744 338014 320896 338042
rect 321020 338014 321172 338042
rect 321296 338014 321448 338042
rect 318950 337742 319024 337770
rect 318892 336728 318944 336734
rect 318892 336670 318944 336676
rect 318524 330472 318576 330478
rect 318524 330414 318576 330420
rect 318904 9042 318932 336670
rect 318996 11762 319024 337742
rect 319088 336734 319116 338014
rect 319076 336728 319128 336734
rect 319076 336670 319128 336676
rect 319364 336122 319392 338014
rect 319352 336116 319404 336122
rect 319352 336058 319404 336064
rect 319076 326936 319128 326942
rect 319076 326878 319128 326884
rect 319088 18698 319116 326878
rect 319640 316034 319668 338014
rect 319916 326942 319944 338014
rect 320192 336258 320220 338014
rect 320468 336666 320496 338014
rect 320456 336660 320508 336666
rect 320456 336602 320508 336608
rect 320180 336252 320232 336258
rect 320180 336194 320232 336200
rect 320744 335354 320772 338014
rect 320824 336116 320876 336122
rect 320824 336058 320876 336064
rect 320376 335326 320772 335354
rect 319904 326936 319956 326942
rect 319904 326878 319956 326884
rect 320272 326596 320324 326602
rect 320272 326538 320324 326544
rect 319180 316006 319668 316034
rect 319076 18692 319128 18698
rect 319076 18634 319128 18640
rect 318984 11756 319036 11762
rect 318984 11698 319036 11704
rect 318892 9036 318944 9042
rect 318892 8978 318944 8984
rect 319180 7614 319208 316006
rect 320284 11830 320312 326538
rect 320376 14618 320404 335326
rect 320456 328092 320508 328098
rect 320456 328034 320508 328040
rect 320364 14612 320416 14618
rect 320364 14554 320416 14560
rect 320272 11824 320324 11830
rect 320272 11766 320324 11772
rect 320468 10334 320496 328034
rect 320456 10328 320508 10334
rect 320456 10270 320508 10276
rect 319168 7608 319220 7614
rect 319168 7550 319220 7556
rect 318524 6180 318576 6186
rect 318524 6122 318576 6128
rect 318064 4888 318116 4894
rect 318064 4830 318116 4836
rect 317328 4208 317380 4214
rect 317328 4150 317380 4156
rect 316224 4072 316276 4078
rect 316224 4014 316276 4020
rect 316236 480 316264 4014
rect 317340 480 317368 4150
rect 318536 480 318564 6122
rect 320836 5030 320864 336058
rect 321020 326602 321048 338014
rect 321296 328098 321324 338014
rect 321710 337770 321738 338028
rect 321848 338014 322000 338042
rect 322124 338014 322276 338042
rect 322400 338014 322552 338042
rect 322676 338014 322828 338042
rect 322952 338014 323104 338042
rect 323228 338014 323380 338042
rect 323504 338014 323656 338042
rect 323780 338014 323932 338042
rect 324056 338014 324208 338042
rect 324332 338014 324484 338042
rect 324608 338014 324760 338042
rect 324884 338014 325036 338042
rect 325160 338014 325312 338042
rect 325436 338014 325588 338042
rect 325804 338014 325864 338042
rect 325988 338014 326140 338042
rect 326264 338014 326416 338042
rect 326540 338014 326692 338042
rect 326816 338014 326968 338042
rect 327244 338014 327396 338042
rect 321710 337742 321784 337770
rect 321652 330540 321704 330546
rect 321652 330482 321704 330488
rect 321284 328092 321336 328098
rect 321284 328034 321336 328040
rect 321008 326596 321060 326602
rect 321008 326538 321060 326544
rect 321664 10402 321692 330482
rect 321652 10396 321704 10402
rect 321652 10338 321704 10344
rect 320916 8968 320968 8974
rect 320916 8910 320968 8916
rect 320824 5024 320876 5030
rect 320824 4966 320876 4972
rect 319720 4140 319772 4146
rect 319720 4082 319772 4088
rect 319732 480 319760 4082
rect 320928 480 320956 8910
rect 321756 7682 321784 337742
rect 321848 336190 321876 338014
rect 322124 336598 322152 338014
rect 322112 336592 322164 336598
rect 322112 336534 322164 336540
rect 322204 336252 322256 336258
rect 322204 336194 322256 336200
rect 321836 336184 321888 336190
rect 321836 336126 321888 336132
rect 321744 7676 321796 7682
rect 321744 7618 321796 7624
rect 322216 4214 322244 336194
rect 322400 330546 322428 338014
rect 322676 336326 322704 338014
rect 322952 336530 322980 338014
rect 322940 336524 322992 336530
rect 322940 336466 322992 336472
rect 322664 336320 322716 336326
rect 322664 336262 322716 336268
rect 323228 335354 323256 338014
rect 323504 336394 323532 338014
rect 323584 336524 323636 336530
rect 323584 336466 323636 336472
rect 323492 336388 323544 336394
rect 323492 336330 323544 336336
rect 323044 335326 323256 335354
rect 322388 330540 322440 330546
rect 322388 330482 322440 330488
rect 322204 4208 322256 4214
rect 322204 4150 322256 4156
rect 323044 3466 323072 335326
rect 323216 330540 323268 330546
rect 323216 330482 323268 330488
rect 323124 329792 323176 329798
rect 323124 329734 323176 329740
rect 323136 51746 323164 329734
rect 323124 51740 323176 51746
rect 323124 51682 323176 51688
rect 323032 3460 323084 3466
rect 323032 3402 323084 3408
rect 322112 3392 322164 3398
rect 322112 3334 322164 3340
rect 322124 480 322152 3334
rect 323228 3330 323256 330482
rect 323596 4962 323624 336466
rect 323676 335436 323728 335442
rect 323676 335378 323728 335384
rect 323688 18630 323716 335378
rect 323780 329798 323808 338014
rect 324056 330546 324084 338014
rect 324332 336054 324360 338014
rect 324608 336530 324636 338014
rect 324596 336524 324648 336530
rect 324596 336466 324648 336472
rect 324320 336048 324372 336054
rect 324320 335990 324372 335996
rect 324044 330540 324096 330546
rect 324044 330482 324096 330488
rect 324412 330540 324464 330546
rect 324412 330482 324464 330488
rect 323768 329792 323820 329798
rect 323768 329734 323820 329740
rect 323676 18624 323728 18630
rect 323676 18566 323728 18572
rect 324424 7818 324452 330482
rect 324504 330472 324556 330478
rect 324504 330414 324556 330420
rect 324516 22778 324544 330414
rect 324884 316034 324912 338014
rect 324964 335368 325016 335374
rect 324964 335310 325016 335316
rect 324608 316006 324912 316034
rect 324504 22772 324556 22778
rect 324504 22714 324556 22720
rect 324412 7812 324464 7818
rect 324412 7754 324464 7760
rect 324412 7608 324464 7614
rect 324412 7550 324464 7556
rect 323584 4956 323636 4962
rect 323584 4898 323636 4904
rect 323308 3596 323360 3602
rect 323308 3538 323360 3544
rect 323216 3324 323268 3330
rect 323216 3266 323268 3272
rect 323320 480 323348 3538
rect 324424 480 324452 7550
rect 324608 3534 324636 316006
rect 324976 17270 325004 335310
rect 325160 330546 325188 338014
rect 325148 330540 325200 330546
rect 325148 330482 325200 330488
rect 325436 330478 325464 338014
rect 325424 330472 325476 330478
rect 325424 330414 325476 330420
rect 324964 17264 325016 17270
rect 324964 17206 325016 17212
rect 325804 3670 325832 338014
rect 325988 335374 326016 338014
rect 325976 335368 326028 335374
rect 326264 335354 326292 338014
rect 325976 335310 326028 335316
rect 326080 335326 326292 335354
rect 326080 330562 326108 335326
rect 325896 330534 326108 330562
rect 325896 294642 325924 330534
rect 326540 316034 326568 338014
rect 326816 335442 326844 338014
rect 326804 335436 326856 335442
rect 326804 335378 326856 335384
rect 327368 330954 327396 338014
rect 327460 338014 327520 338042
rect 327644 338014 327796 338042
rect 327920 338014 328072 338042
rect 328196 338014 328348 338042
rect 327356 330948 327408 330954
rect 327356 330890 327408 330896
rect 327460 330834 327488 338014
rect 327644 335354 327672 338014
rect 327724 336728 327776 336734
rect 327724 336670 327776 336676
rect 325988 316006 326568 316034
rect 327092 330806 327488 330834
rect 327552 335326 327672 335354
rect 325884 294636 325936 294642
rect 325884 294578 325936 294584
rect 325988 3738 326016 316006
rect 327092 3806 327120 330806
rect 327552 330698 327580 335326
rect 327276 330670 327580 330698
rect 327172 330540 327224 330546
rect 327172 330482 327224 330488
rect 327184 3874 327212 330482
rect 327276 13122 327304 330670
rect 327356 330608 327408 330614
rect 327356 330550 327408 330556
rect 327368 292058 327396 330550
rect 327448 330472 327500 330478
rect 327448 330414 327500 330420
rect 327460 318102 327488 330414
rect 327448 318096 327500 318102
rect 327448 318038 327500 318044
rect 327356 292052 327408 292058
rect 327356 291994 327408 292000
rect 327264 13116 327316 13122
rect 327264 13058 327316 13064
rect 327736 6186 327764 336670
rect 327920 330478 327948 338014
rect 328196 330546 328224 338014
rect 328610 337770 328638 338028
rect 328840 338014 328900 338042
rect 329024 338014 329176 338042
rect 329300 338014 329452 338042
rect 329576 338014 329728 338042
rect 329944 338014 330004 338042
rect 330128 338014 330280 338042
rect 330404 338014 330556 338042
rect 330680 338014 330832 338042
rect 330956 338014 331108 338042
rect 331232 338014 331384 338042
rect 331508 338014 331660 338042
rect 331784 338014 331936 338042
rect 332060 338014 332212 338042
rect 332336 338014 332488 338042
rect 332764 338014 332916 338042
rect 328610 337742 328684 337770
rect 328184 330540 328236 330546
rect 328184 330482 328236 330488
rect 327908 330472 327960 330478
rect 327908 330414 327960 330420
rect 328460 330472 328512 330478
rect 328460 330414 328512 330420
rect 327724 6180 327776 6186
rect 327724 6122 327776 6128
rect 328472 3942 328500 330414
rect 328552 325916 328604 325922
rect 328552 325858 328604 325864
rect 328564 10538 328592 325858
rect 328656 14482 328684 337742
rect 328736 330540 328788 330546
rect 328736 330482 328788 330488
rect 328748 21418 328776 330482
rect 328840 285190 328868 338014
rect 329024 330478 329052 338014
rect 329012 330472 329064 330478
rect 329012 330414 329064 330420
rect 329300 325922 329328 338014
rect 329576 330546 329604 338014
rect 329564 330540 329616 330546
rect 329564 330482 329616 330488
rect 329288 325916 329340 325922
rect 329288 325858 329340 325864
rect 328828 285184 328880 285190
rect 328828 285126 328880 285132
rect 328736 21412 328788 21418
rect 328736 21354 328788 21360
rect 328644 14476 328696 14482
rect 328644 14418 328696 14424
rect 328552 10532 328604 10538
rect 328552 10474 328604 10480
rect 329944 4010 329972 338014
rect 330128 336122 330156 338014
rect 330116 336116 330168 336122
rect 330116 336058 330168 336064
rect 330404 335354 330432 338014
rect 330036 335326 330432 335354
rect 330036 278254 330064 335326
rect 330680 316034 330708 338014
rect 330956 336258 330984 338014
rect 331232 336734 331260 338014
rect 331220 336728 331272 336734
rect 331508 336682 331536 338014
rect 331220 336670 331272 336676
rect 331416 336654 331536 336682
rect 330944 336252 330996 336258
rect 330944 336194 330996 336200
rect 331312 330540 331364 330546
rect 331312 330482 331364 330488
rect 330128 316006 330708 316034
rect 330024 278248 330076 278254
rect 330024 278190 330076 278196
rect 330128 4078 330156 316006
rect 330116 4072 330168 4078
rect 330116 4014 330168 4020
rect 329932 4004 329984 4010
rect 329932 3946 329984 3952
rect 328460 3936 328512 3942
rect 328460 3878 328512 3884
rect 327172 3868 327224 3874
rect 327172 3810 327224 3816
rect 327080 3800 327132 3806
rect 327080 3742 327132 3748
rect 328000 3800 328052 3806
rect 328000 3742 328052 3748
rect 325976 3732 326028 3738
rect 325976 3674 326028 3680
rect 325792 3664 325844 3670
rect 325792 3606 325844 3612
rect 324596 3528 324648 3534
rect 324596 3470 324648 3476
rect 326804 3528 326856 3534
rect 326804 3470 326856 3476
rect 325608 3460 325660 3466
rect 325608 3402 325660 3408
rect 325620 480 325648 3402
rect 326816 480 326844 3470
rect 328012 480 328040 3742
rect 331324 3602 331352 330482
rect 331416 4146 331444 336654
rect 331784 335354 331812 338014
rect 331508 335326 331812 335354
rect 331508 8974 331536 335326
rect 332060 316034 332088 338014
rect 332336 330546 332364 338014
rect 332888 335306 332916 338014
rect 332980 338014 333040 338042
rect 333164 338014 333316 338042
rect 333440 338014 333592 338042
rect 333716 338014 333868 338042
rect 334144 338014 334296 338042
rect 332876 335300 332928 335306
rect 332876 335242 332928 335248
rect 332980 330834 333008 338014
rect 333060 335300 333112 335306
rect 333060 335242 333112 335248
rect 332612 330806 333008 330834
rect 332324 330540 332376 330546
rect 332324 330482 332376 330488
rect 331600 316006 332088 316034
rect 331496 8968 331548 8974
rect 331496 8910 331548 8916
rect 331600 6914 331628 316006
rect 331508 6886 331628 6914
rect 331404 4140 331456 4146
rect 331404 4082 331456 4088
rect 331312 3596 331364 3602
rect 331312 3538 331364 3544
rect 331508 3398 331536 6886
rect 331588 3732 331640 3738
rect 331588 3674 331640 3680
rect 331496 3392 331548 3398
rect 331496 3334 331548 3340
rect 329196 3256 329248 3262
rect 329196 3198 329248 3204
rect 329208 480 329236 3198
rect 330392 3188 330444 3194
rect 330392 3130 330444 3136
rect 330404 480 330432 3130
rect 331600 480 331628 3674
rect 332612 3466 332640 330806
rect 332692 330540 332744 330546
rect 332692 330482 332744 330488
rect 332704 3806 332732 330482
rect 332876 330472 332928 330478
rect 332876 330414 332928 330420
rect 332784 330200 332836 330206
rect 332784 330142 332836 330148
rect 332692 3800 332744 3806
rect 332692 3742 332744 3748
rect 332692 3664 332744 3670
rect 332692 3606 332744 3612
rect 332600 3460 332652 3466
rect 332600 3402 332652 3408
rect 332704 480 332732 3606
rect 332796 3262 332824 330142
rect 332888 3534 332916 330414
rect 333072 316034 333100 335242
rect 333164 330478 333192 338014
rect 333440 330546 333468 338014
rect 333428 330540 333480 330546
rect 333428 330482 333480 330488
rect 333152 330472 333204 330478
rect 333152 330414 333204 330420
rect 333716 330206 333744 338014
rect 334072 336728 334124 336734
rect 334072 336670 334124 336676
rect 333980 330472 334032 330478
rect 333980 330414 334032 330420
rect 333704 330200 333756 330206
rect 333704 330142 333756 330148
rect 332980 316006 333100 316034
rect 332980 7614 333008 316006
rect 332968 7608 333020 7614
rect 332968 7550 333020 7556
rect 333992 3602 334020 330414
rect 334084 3738 334112 336670
rect 334268 335354 334296 338014
rect 334360 338014 334420 338042
rect 334544 338014 334696 338042
rect 334820 338014 334972 338042
rect 335096 338014 335248 338042
rect 335372 338014 335524 338042
rect 335648 338014 335800 338042
rect 335924 338014 336076 338042
rect 336200 338014 336352 338042
rect 336476 338014 336628 338042
rect 336904 338014 337056 338042
rect 334360 336734 334388 338014
rect 334348 336728 334400 336734
rect 334348 336670 334400 336676
rect 334544 335354 334572 338014
rect 334268 335326 334388 335354
rect 334360 330818 334388 335326
rect 334452 335326 334572 335354
rect 334348 330812 334400 330818
rect 334348 330754 334400 330760
rect 334452 330698 334480 335326
rect 334176 330670 334480 330698
rect 334072 3732 334124 3738
rect 334072 3674 334124 3680
rect 334176 3670 334204 330670
rect 334348 330608 334400 330614
rect 334348 330550 334400 330556
rect 334256 330540 334308 330546
rect 334256 330482 334308 330488
rect 334164 3664 334216 3670
rect 334164 3606 334216 3612
rect 333980 3596 334032 3602
rect 333980 3538 334032 3544
rect 332876 3528 332928 3534
rect 334268 3482 334296 330482
rect 332876 3470 332928 3476
rect 333900 3454 334296 3482
rect 332784 3256 332836 3262
rect 332784 3198 332836 3204
rect 333900 480 333928 3454
rect 334360 3194 334388 330550
rect 334820 330546 334848 338014
rect 334808 330540 334860 330546
rect 334808 330482 334860 330488
rect 335096 330478 335124 338014
rect 335084 330472 335136 330478
rect 335084 330414 335136 330420
rect 334716 3596 334768 3602
rect 334716 3538 334768 3544
rect 334348 3188 334400 3194
rect 334348 3130 334400 3136
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334728 354 334756 3538
rect 335372 3482 335400 338014
rect 335648 336682 335676 338014
rect 335556 336654 335676 336682
rect 335452 330540 335504 330546
rect 335452 330482 335504 330488
rect 335464 3806 335492 330482
rect 335452 3800 335504 3806
rect 335452 3742 335504 3748
rect 335556 3602 335584 336654
rect 335924 335354 335952 338014
rect 335648 335326 335952 335354
rect 335648 3670 335676 335326
rect 336200 316034 336228 338014
rect 336476 330546 336504 338014
rect 336740 336728 336792 336734
rect 336740 336670 336792 336676
rect 336464 330540 336516 330546
rect 336464 330482 336516 330488
rect 335740 316006 336228 316034
rect 335740 3738 335768 316006
rect 335728 3732 335780 3738
rect 335728 3674 335780 3680
rect 335636 3664 335688 3670
rect 335636 3606 335688 3612
rect 335544 3596 335596 3602
rect 335544 3538 335596 3544
rect 335372 3454 336320 3482
rect 336292 480 336320 3454
rect 336752 2990 336780 336670
rect 336832 330540 336884 330546
rect 336832 330482 336884 330488
rect 336844 3058 336872 330482
rect 336924 330472 336976 330478
rect 336924 330414 336976 330420
rect 336936 4962 336964 330414
rect 336924 4956 336976 4962
rect 336924 4898 336976 4904
rect 337028 4214 337056 338014
rect 337120 338014 337180 338042
rect 337304 338014 337456 338042
rect 337580 338014 337732 338042
rect 337856 338014 338008 338042
rect 338132 338014 338284 338042
rect 338408 338014 338560 338042
rect 338684 338014 338836 338042
rect 338960 338014 339112 338042
rect 339236 338014 339388 338042
rect 337120 336734 337148 338014
rect 337108 336728 337160 336734
rect 337108 336670 337160 336676
rect 337304 330546 337332 338014
rect 337292 330540 337344 330546
rect 337292 330482 337344 330488
rect 337580 330478 337608 338014
rect 337568 330472 337620 330478
rect 337568 330414 337620 330420
rect 337856 316034 337884 338014
rect 337120 316006 337884 316034
rect 337120 21418 337148 316006
rect 337108 21412 337160 21418
rect 337108 21354 337160 21360
rect 337016 4208 337068 4214
rect 337016 4150 337068 4156
rect 337476 3596 337528 3602
rect 337476 3538 337528 3544
rect 336832 3052 336884 3058
rect 336832 2994 336884 3000
rect 336740 2984 336792 2990
rect 336740 2926 336792 2932
rect 337488 480 337516 3538
rect 338132 3534 338160 338014
rect 338212 330540 338264 330546
rect 338212 330482 338264 330488
rect 338120 3528 338172 3534
rect 338120 3470 338172 3476
rect 338224 3466 338252 330482
rect 338304 330472 338356 330478
rect 338304 330414 338356 330420
rect 338316 4894 338344 330414
rect 338408 7682 338436 338014
rect 338684 316742 338712 338014
rect 338960 330546 338988 338014
rect 338948 330540 339000 330546
rect 338948 330482 339000 330488
rect 339236 330478 339264 338014
rect 339650 337770 339678 338028
rect 339940 338014 340092 338042
rect 339650 337742 339724 337770
rect 339500 330540 339552 330546
rect 339500 330482 339552 330488
rect 339224 330472 339276 330478
rect 339224 330414 339276 330420
rect 338672 316736 338724 316742
rect 338672 316678 338724 316684
rect 338396 7676 338448 7682
rect 338396 7618 338448 7624
rect 339512 6186 339540 330482
rect 339592 328092 339644 328098
rect 339592 328034 339644 328040
rect 339604 14482 339632 328034
rect 339696 305658 339724 337742
rect 340064 336326 340092 338014
rect 340156 338014 340216 338042
rect 340340 338014 340492 338042
rect 340616 338014 340768 338042
rect 340892 338014 341044 338042
rect 341260 338014 341320 338042
rect 341444 338014 341596 338042
rect 341720 338014 341872 338042
rect 342088 338014 342148 338042
rect 342364 338014 342424 338042
rect 342548 338014 342700 338042
rect 342824 338014 342976 338042
rect 343100 338014 343252 338042
rect 343376 338014 343528 338042
rect 343744 338014 343804 338042
rect 343928 338014 344080 338042
rect 344296 338014 344356 338042
rect 344480 338014 344632 338042
rect 344756 338014 344908 338042
rect 345124 338014 345184 338042
rect 345308 338014 345460 338042
rect 345584 338014 345736 338042
rect 345860 338014 346012 338042
rect 346136 338014 346288 338042
rect 346564 338014 346716 338042
rect 340052 336320 340104 336326
rect 340052 336262 340104 336268
rect 340156 336258 340184 338014
rect 340144 336252 340196 336258
rect 340144 336194 340196 336200
rect 340340 328098 340368 338014
rect 340616 330546 340644 338014
rect 340604 330540 340656 330546
rect 340604 330482 340656 330488
rect 340328 328092 340380 328098
rect 340328 328034 340380 328040
rect 339684 305652 339736 305658
rect 339684 305594 339736 305600
rect 339592 14476 339644 14482
rect 339592 14418 339644 14424
rect 340892 8974 340920 338014
rect 341260 336054 341288 338014
rect 341248 336048 341300 336054
rect 341248 335990 341300 335996
rect 340972 326392 341024 326398
rect 340972 326334 341024 326340
rect 340984 11762 341012 326334
rect 341444 316034 341472 338014
rect 341524 336320 341576 336326
rect 341524 336262 341576 336268
rect 341076 316006 341472 316034
rect 341076 24138 341104 316006
rect 341536 269822 341564 336262
rect 341720 326398 341748 338014
rect 342088 336462 342116 338014
rect 342076 336456 342128 336462
rect 342076 336398 342128 336404
rect 342364 336122 342392 338014
rect 342352 336116 342404 336122
rect 342352 336058 342404 336064
rect 342548 335354 342576 338014
rect 342272 335326 342576 335354
rect 341708 326392 341760 326398
rect 341708 326334 341760 326340
rect 341524 269816 341576 269822
rect 341524 269758 341576 269764
rect 341064 24132 341116 24138
rect 341064 24074 341116 24080
rect 340972 11756 341024 11762
rect 340972 11698 341024 11704
rect 340880 8968 340932 8974
rect 340880 8910 340932 8916
rect 339500 6180 339552 6186
rect 339500 6122 339552 6128
rect 338304 4888 338356 4894
rect 338304 4830 338356 4836
rect 342272 4826 342300 335326
rect 342352 326392 342404 326398
rect 342352 326334 342404 326340
rect 342364 10334 342392 326334
rect 342444 323604 342496 323610
rect 342444 323546 342496 323552
rect 342456 22778 342484 323546
rect 342824 316034 342852 338014
rect 343100 323610 343128 338014
rect 343376 326398 343404 338014
rect 343744 335850 343772 338014
rect 343732 335844 343784 335850
rect 343732 335786 343784 335792
rect 343364 326392 343416 326398
rect 343364 326334 343416 326340
rect 343640 326392 343692 326398
rect 343640 326334 343692 326340
rect 343088 323604 343140 323610
rect 343088 323546 343140 323552
rect 342548 316006 342852 316034
rect 342548 291854 342576 316006
rect 342536 291848 342588 291854
rect 342536 291790 342588 291796
rect 343652 25566 343680 326334
rect 343732 324420 343784 324426
rect 343732 324362 343784 324368
rect 343744 284986 343772 324362
rect 343928 316034 343956 338014
rect 344296 336530 344324 338014
rect 344284 336524 344336 336530
rect 344284 336466 344336 336472
rect 344480 324426 344508 338014
rect 344756 326398 344784 338014
rect 345124 336326 345152 338014
rect 345112 336320 345164 336326
rect 345112 336262 345164 336268
rect 345204 326460 345256 326466
rect 345204 326402 345256 326408
rect 344744 326392 344796 326398
rect 344744 326334 344796 326340
rect 345112 326392 345164 326398
rect 345112 326334 345164 326340
rect 345020 326324 345072 326330
rect 345020 326266 345072 326272
rect 344468 324420 344520 324426
rect 344468 324362 344520 324368
rect 343836 316006 343956 316034
rect 343836 313954 343864 316006
rect 343824 313948 343876 313954
rect 343824 313890 343876 313896
rect 343732 284980 343784 284986
rect 343732 284922 343784 284928
rect 343640 25560 343692 25566
rect 343640 25502 343692 25508
rect 342444 22772 342496 22778
rect 342444 22714 342496 22720
rect 342352 10328 342404 10334
rect 342352 10270 342404 10276
rect 345032 7614 345060 326266
rect 345124 15978 345152 326334
rect 345216 47734 345244 326402
rect 345308 307086 345336 338014
rect 345584 326398 345612 338014
rect 345664 335844 345716 335850
rect 345664 335786 345716 335792
rect 345572 326392 345624 326398
rect 345572 326334 345624 326340
rect 345296 307080 345348 307086
rect 345296 307022 345348 307028
rect 345676 287706 345704 335786
rect 345860 326330 345888 338014
rect 346136 326466 346164 338014
rect 346688 328454 346716 338014
rect 346780 338014 346840 338042
rect 346964 338014 347116 338042
rect 347240 338014 347392 338042
rect 347516 338014 347668 338042
rect 346780 336394 346808 338014
rect 346768 336388 346820 336394
rect 346768 336330 346820 336336
rect 346964 335354 346992 338014
rect 346596 328426 346716 328454
rect 346780 335326 346992 335354
rect 346124 326460 346176 326466
rect 346124 326402 346176 326408
rect 346400 326460 346452 326466
rect 346400 326402 346452 326408
rect 345848 326324 345900 326330
rect 345848 326266 345900 326272
rect 345664 287700 345716 287706
rect 345664 287642 345716 287648
rect 345204 47728 345256 47734
rect 345204 47670 345256 47676
rect 345112 15972 345164 15978
rect 345112 15914 345164 15920
rect 346412 13190 346440 326402
rect 346492 326392 346544 326398
rect 346492 326334 346544 326340
rect 346504 140078 346532 326334
rect 346596 322946 346624 328426
rect 346596 322918 346716 322946
rect 346584 321700 346636 321706
rect 346584 321642 346636 321648
rect 346596 278050 346624 321642
rect 346688 279478 346716 322918
rect 346780 321706 346808 335326
rect 347240 326398 347268 338014
rect 347516 326466 347544 338014
rect 347930 337770 347958 338028
rect 348068 338014 348220 338042
rect 348496 338014 348648 338042
rect 347930 337742 348004 337770
rect 347976 326466 348004 337742
rect 347504 326460 347556 326466
rect 347504 326402 347556 326408
rect 347964 326460 348016 326466
rect 347964 326402 348016 326408
rect 347228 326392 347280 326398
rect 347228 326334 347280 326340
rect 347780 326392 347832 326398
rect 347780 326334 347832 326340
rect 346768 321700 346820 321706
rect 346768 321642 346820 321648
rect 346676 279472 346728 279478
rect 346676 279414 346728 279420
rect 346584 278044 346636 278050
rect 346584 277986 346636 277992
rect 346492 140072 346544 140078
rect 346492 140014 346544 140020
rect 347792 26926 347820 326334
rect 348068 323626 348096 338014
rect 348620 336734 348648 338014
rect 348712 338014 348772 338042
rect 348896 338014 349048 338042
rect 349264 338014 349324 338042
rect 348608 336728 348660 336734
rect 348608 336670 348660 336676
rect 348712 336598 348740 338014
rect 348700 336592 348752 336598
rect 348700 336534 348752 336540
rect 348148 326460 348200 326466
rect 348148 326402 348200 326408
rect 347884 323598 348096 323626
rect 347884 271182 347912 323598
rect 348160 318794 348188 326402
rect 348896 326398 348924 338014
rect 348884 326392 348936 326398
rect 348884 326334 348936 326340
rect 349160 326392 349212 326398
rect 349160 326334 349212 326340
rect 347976 318766 348188 318794
rect 347976 311302 348004 318766
rect 347964 311296 348016 311302
rect 347964 311238 348016 311244
rect 347872 271176 347924 271182
rect 347872 271118 347924 271124
rect 347780 26920 347832 26926
rect 347780 26862 347832 26868
rect 346492 21412 346544 21418
rect 346492 21354 346544 21360
rect 346504 16574 346532 21354
rect 349172 17338 349200 326334
rect 349264 322386 349292 338014
rect 349586 337770 349614 338028
rect 349724 338014 349876 338042
rect 350000 338014 350152 338042
rect 350276 338014 350428 338042
rect 350552 338014 350704 338042
rect 350828 338014 350980 338042
rect 351104 338014 351256 338042
rect 351380 338014 351532 338042
rect 351656 338014 351808 338042
rect 352024 338014 352084 338042
rect 352208 338014 352360 338042
rect 352484 338014 352636 338042
rect 352760 338014 352912 338042
rect 353036 338014 353188 338042
rect 353464 338014 353616 338042
rect 349586 337742 349660 337770
rect 349632 332042 349660 337742
rect 349620 332036 349672 332042
rect 349620 331978 349672 331984
rect 349724 331214 349752 338014
rect 349804 336728 349856 336734
rect 349804 336670 349856 336676
rect 349356 331186 349752 331214
rect 349252 322380 349304 322386
rect 349252 322322 349304 322328
rect 349252 316736 349304 316742
rect 349252 316678 349304 316684
rect 349160 17332 349212 17338
rect 349160 17274 349212 17280
rect 346504 16546 346992 16574
rect 346400 13184 346452 13190
rect 346400 13126 346452 13132
rect 345020 7608 345072 7614
rect 345020 7550 345072 7556
rect 345756 4956 345808 4962
rect 345756 4898 345808 4904
rect 342260 4820 342312 4826
rect 342260 4762 342312 4768
rect 342168 4208 342220 4214
rect 342168 4150 342220 4156
rect 340972 3800 341024 3806
rect 340972 3742 341024 3748
rect 339868 3732 339920 3738
rect 339868 3674 339920 3680
rect 338672 3664 338724 3670
rect 338672 3606 338724 3612
rect 338212 3460 338264 3466
rect 338212 3402 338264 3408
rect 338684 480 338712 3606
rect 339880 480 339908 3674
rect 340984 480 341012 3742
rect 342180 480 342208 4150
rect 344560 3052 344612 3058
rect 344560 2994 344612 3000
rect 343364 2984 343416 2990
rect 343364 2926 343416 2932
rect 343376 480 343404 2926
rect 344572 480 344600 2994
rect 345768 480 345796 4898
rect 346964 480 346992 16546
rect 349160 7676 349212 7682
rect 349160 7618 349212 7624
rect 348056 3528 348108 3534
rect 348056 3470 348108 3476
rect 348068 480 348096 3470
rect 349172 3346 349200 7618
rect 349264 3534 349292 316678
rect 349356 28286 349384 331186
rect 349816 325106 349844 336670
rect 349804 325100 349856 325106
rect 349804 325042 349856 325048
rect 350000 321554 350028 338014
rect 350276 326398 350304 338014
rect 350264 326392 350316 326398
rect 350264 326334 350316 326340
rect 349448 321526 350028 321554
rect 349448 316878 349476 321526
rect 349436 316872 349488 316878
rect 349436 316814 349488 316820
rect 350552 86290 350580 338014
rect 350724 326460 350776 326466
rect 350724 326402 350776 326408
rect 350632 326392 350684 326398
rect 350632 326334 350684 326340
rect 350644 178702 350672 326334
rect 350736 309942 350764 326402
rect 350828 326346 350856 338014
rect 351104 335354 351132 338014
rect 351012 335326 351132 335354
rect 351012 326466 351040 335326
rect 351000 326460 351052 326466
rect 351000 326402 351052 326408
rect 351380 326398 351408 338014
rect 351368 326392 351420 326398
rect 350828 326318 350948 326346
rect 351368 326334 351420 326340
rect 350816 326256 350868 326262
rect 350816 326198 350868 326204
rect 350828 319598 350856 326198
rect 350920 321026 350948 326318
rect 351656 326262 351684 338014
rect 352024 330682 352052 338014
rect 352208 335354 352236 338014
rect 352116 335326 352236 335354
rect 352012 330676 352064 330682
rect 352012 330618 352064 330624
rect 351920 326392 351972 326398
rect 352116 326380 352144 335326
rect 351920 326334 351972 326340
rect 352024 326352 352144 326380
rect 351644 326256 351696 326262
rect 351644 326198 351696 326204
rect 350908 321020 350960 321026
rect 350908 320962 350960 320968
rect 350816 319592 350868 319598
rect 350816 319534 350868 319540
rect 350724 309936 350776 309942
rect 350724 309878 350776 309884
rect 350632 178696 350684 178702
rect 350632 178638 350684 178644
rect 350540 86284 350592 86290
rect 350540 86226 350592 86232
rect 349344 28280 349396 28286
rect 349344 28222 349396 28228
rect 351932 11830 351960 326334
rect 352024 29646 352052 326352
rect 352484 325038 352512 338014
rect 352472 325032 352524 325038
rect 352472 324974 352524 324980
rect 352760 321554 352788 338014
rect 353036 326398 353064 338014
rect 353484 336728 353536 336734
rect 353484 336670 353536 336676
rect 353392 326460 353444 326466
rect 353392 326402 353444 326408
rect 353024 326392 353076 326398
rect 353024 326334 353076 326340
rect 353300 326392 353352 326398
rect 353300 326334 353352 326340
rect 352116 321526 352788 321554
rect 352116 308514 352144 321526
rect 352104 308508 352156 308514
rect 352104 308450 352156 308456
rect 352012 29640 352064 29646
rect 352012 29582 352064 29588
rect 351920 11824 351972 11830
rect 351920 11766 351972 11772
rect 353312 4894 353340 326334
rect 353404 312594 353432 326402
rect 353392 312588 353444 312594
rect 353392 312530 353444 312536
rect 353392 305652 353444 305658
rect 353392 305594 353444 305600
rect 353404 16574 353432 305594
rect 353496 272542 353524 336670
rect 353588 335354 353616 338014
rect 353680 338014 353740 338042
rect 353864 338014 354016 338042
rect 354140 338014 354292 338042
rect 354416 338014 354568 338042
rect 353680 336734 353708 338014
rect 353668 336728 353720 336734
rect 353668 336670 353720 336676
rect 353588 335326 353708 335354
rect 353680 323746 353708 335326
rect 353864 326398 353892 338014
rect 353852 326392 353904 326398
rect 353852 326334 353904 326340
rect 353668 323740 353720 323746
rect 353668 323682 353720 323688
rect 354140 321554 354168 338014
rect 354416 326466 354444 338014
rect 354830 337770 354858 338028
rect 355060 338014 355120 338042
rect 355244 338014 355396 338042
rect 355520 338014 355672 338042
rect 355796 338014 355948 338042
rect 356224 338014 356376 338042
rect 354830 337742 354904 337770
rect 354404 326460 354456 326466
rect 354404 326402 354456 326408
rect 354772 326460 354824 326466
rect 354772 326402 354824 326408
rect 354680 322788 354732 322794
rect 354680 322730 354732 322736
rect 353588 321526 354168 321554
rect 353588 305794 353616 321526
rect 353576 305788 353628 305794
rect 353576 305730 353628 305736
rect 354692 304366 354720 322730
rect 354680 304360 354732 304366
rect 354680 304302 354732 304308
rect 353484 272536 353536 272542
rect 353484 272478 353536 272484
rect 354680 269816 354732 269822
rect 354680 269758 354732 269764
rect 354692 16574 354720 269758
rect 354784 244934 354812 326402
rect 354876 258738 354904 337742
rect 354956 326392 355008 326398
rect 354956 326334 355008 326340
rect 354968 269890 354996 326334
rect 355060 318238 355088 338014
rect 355244 326398 355272 338014
rect 355520 326466 355548 338014
rect 355508 326460 355560 326466
rect 355508 326402 355560 326408
rect 355232 326392 355284 326398
rect 355232 326334 355284 326340
rect 355796 322794 355824 338014
rect 356244 336728 356296 336734
rect 356244 336670 356296 336676
rect 356060 336252 356112 336258
rect 356060 336194 356112 336200
rect 355784 322788 355836 322794
rect 355784 322730 355836 322736
rect 355048 318232 355100 318238
rect 355048 318174 355100 318180
rect 354956 269884 355008 269890
rect 354956 269826 355008 269832
rect 354864 258732 354916 258738
rect 354864 258674 354916 258680
rect 354772 244928 354824 244934
rect 354772 244870 354824 244876
rect 353404 16546 353616 16574
rect 354692 16546 355272 16574
rect 352840 4888 352892 4894
rect 352840 4830 352892 4836
rect 353300 4888 353352 4894
rect 353300 4830 353352 4836
rect 349252 3528 349304 3534
rect 349252 3470 349304 3476
rect 350448 3528 350500 3534
rect 350448 3470 350500 3476
rect 349172 3318 349292 3346
rect 349264 480 349292 3318
rect 350460 480 350488 3470
rect 351644 3460 351696 3466
rect 351644 3402 351696 3408
rect 351656 480 351684 3402
rect 352852 480 352880 4830
rect 335054 354 335166 480
rect 334728 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 353588 354 353616 16546
rect 355244 480 355272 16546
rect 356072 3482 356100 336194
rect 356152 326392 356204 326398
rect 356152 326334 356204 326340
rect 356164 3602 356192 326334
rect 356256 16574 356284 336670
rect 356348 335354 356376 338014
rect 356440 338014 356500 338042
rect 356716 338014 356776 338042
rect 356900 338014 357052 338042
rect 357176 338014 357328 338042
rect 357544 338014 357604 338042
rect 357728 338014 357880 338042
rect 358004 338014 358156 338042
rect 358280 338014 358432 338042
rect 358556 338014 358708 338042
rect 358924 338014 358984 338042
rect 359108 338014 359260 338042
rect 359384 338014 359536 338042
rect 359660 338014 359812 338042
rect 359936 338014 360088 338042
rect 360364 338014 360516 338042
rect 356440 336734 356468 338014
rect 356428 336728 356480 336734
rect 356428 336670 356480 336676
rect 356716 335918 356744 338014
rect 356704 335912 356756 335918
rect 356704 335854 356756 335860
rect 356348 335326 356468 335354
rect 356336 323196 356388 323202
rect 356336 323138 356388 323144
rect 356348 307154 356376 323138
rect 356440 316810 356468 335326
rect 356900 323202 356928 338014
rect 357176 326398 357204 338014
rect 357544 335782 357572 338014
rect 357532 335776 357584 335782
rect 357532 335718 357584 335724
rect 357532 326460 357584 326466
rect 357532 326402 357584 326408
rect 357164 326392 357216 326398
rect 357164 326334 357216 326340
rect 357440 326392 357492 326398
rect 357440 326334 357492 326340
rect 356888 323196 356940 323202
rect 356888 323138 356940 323144
rect 356428 316804 356480 316810
rect 356428 316746 356480 316752
rect 356336 307148 356388 307154
rect 356336 307090 356388 307096
rect 356256 16546 356468 16574
rect 356152 3596 356204 3602
rect 356152 3538 356204 3544
rect 356072 3454 356376 3482
rect 356348 480 356376 3454
rect 356440 3262 356468 16546
rect 357452 3398 357480 326334
rect 357544 303006 357572 326402
rect 357624 326324 357676 326330
rect 357624 326266 357676 326272
rect 357636 311234 357664 326266
rect 357728 319530 357756 338014
rect 358004 326398 358032 338014
rect 358280 326466 358308 338014
rect 358268 326460 358320 326466
rect 358268 326402 358320 326408
rect 357992 326392 358044 326398
rect 357992 326334 358044 326340
rect 358556 326330 358584 338014
rect 358924 336258 358952 338014
rect 358912 336252 358964 336258
rect 358912 336194 358964 336200
rect 358912 326460 358964 326466
rect 358912 326402 358964 326408
rect 358820 326392 358872 326398
rect 358820 326334 358872 326340
rect 358544 326324 358596 326330
rect 358544 326266 358596 326272
rect 357716 319524 357768 319530
rect 357716 319466 357768 319472
rect 357624 311228 357676 311234
rect 357624 311170 357676 311176
rect 357532 303000 357584 303006
rect 357532 302942 357584 302948
rect 357532 14476 357584 14482
rect 357532 14418 357584 14424
rect 357440 3392 357492 3398
rect 357440 3334 357492 3340
rect 356428 3256 356480 3262
rect 356428 3198 356480 3204
rect 357544 480 357572 14418
rect 358728 6180 358780 6186
rect 358728 6122 358780 6128
rect 358740 480 358768 6122
rect 358832 4146 358860 326334
rect 358924 300218 358952 326402
rect 359108 316034 359136 338014
rect 359384 334762 359412 338014
rect 359556 336524 359608 336530
rect 359556 336466 359608 336472
rect 359464 336048 359516 336054
rect 359464 335990 359516 335996
rect 359372 334756 359424 334762
rect 359372 334698 359424 334704
rect 359016 316006 359136 316034
rect 359016 301578 359044 316006
rect 359004 301572 359056 301578
rect 359004 301514 359056 301520
rect 358912 300212 358964 300218
rect 358912 300154 358964 300160
rect 359476 9654 359504 335990
rect 359568 323610 359596 336466
rect 359660 326398 359688 338014
rect 359936 326466 359964 338014
rect 360488 333402 360516 338014
rect 360580 338014 360640 338042
rect 360764 338014 360916 338042
rect 361040 338014 361192 338042
rect 361316 338014 361468 338042
rect 361684 338014 361744 338042
rect 361868 338014 362020 338042
rect 362236 338014 362296 338042
rect 362420 338014 362572 338042
rect 362696 338014 362848 338042
rect 362972 338014 363124 338042
rect 363248 338014 363400 338042
rect 363524 338014 363676 338042
rect 363892 338014 363952 338042
rect 364076 338014 364228 338042
rect 364504 338014 364656 338042
rect 360580 336190 360608 338014
rect 360568 336184 360620 336190
rect 360568 336126 360620 336132
rect 360568 335912 360620 335918
rect 360568 335854 360620 335860
rect 360476 333396 360528 333402
rect 360476 333338 360528 333344
rect 360292 330540 360344 330546
rect 360292 330482 360344 330488
rect 360200 330472 360252 330478
rect 360200 330414 360252 330420
rect 359924 326460 359976 326466
rect 359924 326402 359976 326408
rect 359648 326392 359700 326398
rect 359648 326334 359700 326340
rect 359556 323604 359608 323610
rect 359556 323546 359608 323552
rect 359464 9648 359516 9654
rect 359464 9590 359516 9596
rect 359924 8968 359976 8974
rect 359924 8910 359976 8916
rect 358820 4140 358872 4146
rect 358820 4082 358872 4088
rect 359936 480 359964 8910
rect 360212 4078 360240 330414
rect 360304 268394 360332 330482
rect 360580 329254 360608 335854
rect 360568 329248 360620 329254
rect 360568 329190 360620 329196
rect 360764 316034 360792 338014
rect 360844 336116 360896 336122
rect 360844 336058 360896 336064
rect 360396 316006 360792 316034
rect 360396 298858 360424 316006
rect 360384 298852 360436 298858
rect 360384 298794 360436 298800
rect 360292 268388 360344 268394
rect 360292 268330 360344 268336
rect 360856 8430 360884 336058
rect 360936 335776 360988 335782
rect 360936 335718 360988 335724
rect 360948 315450 360976 335718
rect 361040 330546 361068 338014
rect 361028 330540 361080 330546
rect 361028 330482 361080 330488
rect 361316 330478 361344 338014
rect 361684 335714 361712 338014
rect 361672 335708 361724 335714
rect 361672 335650 361724 335656
rect 361580 330540 361632 330546
rect 361580 330482 361632 330488
rect 361304 330472 361356 330478
rect 361304 330414 361356 330420
rect 360936 315444 360988 315450
rect 360936 315386 360988 315392
rect 361592 267034 361620 330482
rect 361672 327956 361724 327962
rect 361672 327898 361724 327904
rect 361684 297498 361712 327898
rect 361868 318170 361896 338014
rect 362236 336122 362264 338014
rect 362224 336116 362276 336122
rect 362224 336058 362276 336064
rect 362420 327962 362448 338014
rect 362696 330546 362724 338014
rect 362684 330540 362736 330546
rect 362684 330482 362736 330488
rect 362408 327956 362460 327962
rect 362408 327898 362460 327904
rect 361856 318164 361908 318170
rect 361856 318106 361908 318112
rect 361672 297492 361724 297498
rect 361672 297434 361724 297440
rect 361580 267028 361632 267034
rect 361580 266970 361632 266976
rect 361580 24132 361632 24138
rect 361580 24074 361632 24080
rect 361592 16574 361620 24074
rect 361592 16546 361896 16574
rect 361120 9648 361172 9654
rect 361120 9590 361172 9596
rect 360844 8424 360896 8430
rect 360844 8366 360896 8372
rect 360200 4072 360252 4078
rect 360200 4014 360252 4020
rect 361132 480 361160 9590
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 361868 354 361896 16546
rect 362972 4010 363000 338014
rect 363144 330540 363196 330546
rect 363144 330482 363196 330488
rect 363052 326664 363104 326670
rect 363052 326606 363104 326612
rect 363064 265674 363092 326606
rect 363156 294710 363184 330482
rect 363248 296070 363276 338014
rect 363524 326670 363552 338014
rect 363604 336456 363656 336462
rect 363604 336398 363656 336404
rect 363512 326664 363564 326670
rect 363512 326606 363564 326612
rect 363236 296064 363288 296070
rect 363236 296006 363288 296012
rect 363144 294704 363196 294710
rect 363144 294646 363196 294652
rect 363052 265668 363104 265674
rect 363052 265610 363104 265616
rect 363512 11756 363564 11762
rect 363512 11698 363564 11704
rect 362960 4004 363012 4010
rect 362960 3946 363012 3952
rect 363524 480 363552 11698
rect 363616 4826 363644 336398
rect 363892 336054 363920 338014
rect 363880 336048 363932 336054
rect 363880 335990 363932 335996
rect 363696 335708 363748 335714
rect 363696 335650 363748 335656
rect 363708 327826 363736 335650
rect 364076 330546 364104 338014
rect 364064 330540 364116 330546
rect 364064 330482 364116 330488
rect 364524 330540 364576 330546
rect 364524 330482 364576 330488
rect 364432 330472 364484 330478
rect 364432 330414 364484 330420
rect 364248 328568 364300 328574
rect 364248 328510 364300 328516
rect 364260 328454 364288 328510
rect 364260 328426 364380 328454
rect 363696 327820 363748 327826
rect 363696 327762 363748 327768
rect 363604 4820 363656 4826
rect 363604 4762 363656 4768
rect 364352 3942 364380 328426
rect 364340 3936 364392 3942
rect 364340 3878 364392 3884
rect 364444 3874 364472 330414
rect 364536 264246 364564 330482
rect 364628 309874 364656 338014
rect 364720 338014 364780 338042
rect 364904 338014 365056 338042
rect 365180 338014 365332 338042
rect 365456 338014 365608 338042
rect 365824 338014 365884 338042
rect 366008 338014 366160 338042
rect 366284 338014 366436 338042
rect 366560 338014 366712 338042
rect 366836 338014 366988 338042
rect 367112 338014 367264 338042
rect 367388 338014 367540 338042
rect 367664 338014 367816 338042
rect 367940 338014 368092 338042
rect 368216 338014 368368 338042
rect 364720 328574 364748 338014
rect 364708 328568 364760 328574
rect 364708 328510 364760 328516
rect 364904 326466 364932 338014
rect 365180 330546 365208 338014
rect 365168 330540 365220 330546
rect 365168 330482 365220 330488
rect 365456 330478 365484 338014
rect 365824 335918 365852 338014
rect 365812 335912 365864 335918
rect 365812 335854 365864 335860
rect 366008 335354 366036 338014
rect 365916 335326 366036 335354
rect 365720 330540 365772 330546
rect 365720 330482 365772 330488
rect 365444 330472 365496 330478
rect 365444 330414 365496 330420
rect 364892 326460 364944 326466
rect 364892 326402 364944 326408
rect 364616 309868 364668 309874
rect 364616 309810 364668 309816
rect 364524 264240 364576 264246
rect 364524 264182 364576 264188
rect 364616 4820 364668 4826
rect 364616 4762 364668 4768
rect 364432 3868 364484 3874
rect 364432 3810 364484 3816
rect 364628 480 364656 4762
rect 365732 3806 365760 330482
rect 365812 330472 365864 330478
rect 365812 330414 365864 330420
rect 365824 296002 365852 330414
rect 365916 315382 365944 335326
rect 366284 330546 366312 338014
rect 366272 330540 366324 330546
rect 366272 330482 366324 330488
rect 366560 322318 366588 338014
rect 366836 330478 366864 338014
rect 366824 330472 366876 330478
rect 366824 330414 366876 330420
rect 366548 322312 366600 322318
rect 366548 322254 366600 322260
rect 365904 315376 365956 315382
rect 365904 315318 365956 315324
rect 365812 295996 365864 296002
rect 365812 295938 365864 295944
rect 365812 8424 365864 8430
rect 365812 8366 365864 8372
rect 365720 3800 365772 3806
rect 365720 3742 365772 3748
rect 365824 480 365852 8366
rect 367008 4752 367060 4758
rect 367008 4694 367060 4700
rect 367020 480 367048 4694
rect 367112 3738 367140 338014
rect 367388 336682 367416 338014
rect 367296 336654 367416 336682
rect 367192 328228 367244 328234
rect 367192 328170 367244 328176
rect 367100 3732 367152 3738
rect 367100 3674 367152 3680
rect 367204 3670 367232 328170
rect 367296 305726 367324 336654
rect 367664 335354 367692 338014
rect 367388 335326 367692 335354
rect 367284 305720 367336 305726
rect 367284 305662 367336 305668
rect 367284 291848 367336 291854
rect 367284 291790 367336 291796
rect 367296 16574 367324 291790
rect 367388 262886 367416 335326
rect 367940 328234 367968 338014
rect 367928 328228 367980 328234
rect 367928 328170 367980 328176
rect 368216 316034 368244 338014
rect 368630 337770 368658 338028
rect 368768 338014 368920 338042
rect 368630 337742 368704 337770
rect 368480 330540 368532 330546
rect 368480 330482 368532 330488
rect 367480 316006 368244 316034
rect 367480 291922 367508 316006
rect 367468 291916 367520 291922
rect 367468 291858 367520 291864
rect 367376 262880 367428 262886
rect 367376 262822 367428 262828
rect 367296 16546 367784 16574
rect 367192 3664 367244 3670
rect 367192 3606 367244 3612
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 16546
rect 368492 3534 368520 330482
rect 368572 330472 368624 330478
rect 368572 330414 368624 330420
rect 368584 18630 368612 330414
rect 368676 261526 368704 337742
rect 368768 330546 368796 338014
rect 369182 337770 369210 338028
rect 369320 338014 369472 338042
rect 369596 338014 369748 338042
rect 369964 338014 370024 338042
rect 370148 338014 370300 338042
rect 370424 338014 370576 338042
rect 370792 338014 370852 338042
rect 370976 338014 371128 338042
rect 371252 338014 371404 338042
rect 369182 337742 369256 337770
rect 369124 335912 369176 335918
rect 369124 335854 369176 335860
rect 368756 330540 368808 330546
rect 368756 330482 368808 330488
rect 368756 325916 368808 325922
rect 368756 325858 368808 325864
rect 368768 314022 368796 325858
rect 368756 314016 368808 314022
rect 368756 313958 368808 313964
rect 369136 293350 369164 335854
rect 369228 334694 369256 337742
rect 369216 334688 369268 334694
rect 369216 334630 369268 334636
rect 369320 325922 369348 338014
rect 369596 330478 369624 338014
rect 369964 336462 369992 338014
rect 369952 336456 370004 336462
rect 369952 336398 370004 336404
rect 369584 330472 369636 330478
rect 369584 330414 369636 330420
rect 369860 326392 369912 326398
rect 369860 326334 369912 326340
rect 369308 325916 369360 325922
rect 369308 325858 369360 325864
rect 369124 293344 369176 293350
rect 369124 293286 369176 293292
rect 368664 261520 368716 261526
rect 368664 261462 368716 261468
rect 369872 260166 369900 326334
rect 369952 326324 370004 326330
rect 369952 326266 370004 326272
rect 369964 289134 369992 326266
rect 370148 316034 370176 338014
rect 370424 326398 370452 338014
rect 370504 336592 370556 336598
rect 370504 336534 370556 336540
rect 370412 326392 370464 326398
rect 370412 326334 370464 326340
rect 370056 316006 370176 316034
rect 370056 290562 370084 316006
rect 370044 290556 370096 290562
rect 370044 290498 370096 290504
rect 369952 289128 370004 289134
rect 369952 289070 370004 289076
rect 369860 260160 369912 260166
rect 369860 260102 369912 260108
rect 368664 22772 368716 22778
rect 368664 22714 368716 22720
rect 368572 18624 368624 18630
rect 368572 18566 368624 18572
rect 368676 16574 368704 22714
rect 368676 16546 369440 16574
rect 368480 3528 368532 3534
rect 368480 3470 368532 3476
rect 369412 480 369440 16546
rect 370136 10328 370188 10334
rect 370136 10270 370188 10276
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370148 354 370176 10270
rect 370516 8974 370544 336534
rect 370792 336530 370820 338014
rect 370780 336524 370832 336530
rect 370780 336466 370832 336472
rect 370976 326330 371004 338014
rect 370964 326324 371016 326330
rect 370964 326266 371016 326272
rect 371252 294642 371280 338014
rect 371666 337770 371694 338028
rect 371804 338014 371956 338042
rect 372080 338014 372232 338042
rect 371666 337742 371740 337770
rect 371712 331974 371740 337742
rect 371700 331968 371752 331974
rect 371700 331910 371752 331916
rect 371332 326392 371384 326398
rect 371332 326334 371384 326340
rect 371240 294636 371292 294642
rect 371240 294578 371292 294584
rect 371240 287700 371292 287706
rect 371240 287642 371292 287648
rect 370504 8968 370556 8974
rect 370504 8910 370556 8916
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 371252 354 371280 287642
rect 371344 257378 371372 326334
rect 371804 316034 371832 338014
rect 371884 336320 371936 336326
rect 371884 336262 371936 336268
rect 371436 316006 371832 316034
rect 371436 287706 371464 316006
rect 371424 287700 371476 287706
rect 371424 287642 371476 287648
rect 371332 257372 371384 257378
rect 371332 257314 371384 257320
rect 371896 4826 371924 336262
rect 372080 326398 372108 338014
rect 372494 337770 372522 338028
rect 372784 338014 372936 338042
rect 372494 337742 372568 337770
rect 372540 333130 372568 337742
rect 372712 336728 372764 336734
rect 372712 336670 372764 336676
rect 372528 333124 372580 333130
rect 372528 333066 372580 333072
rect 372068 326392 372120 326398
rect 372068 326334 372120 326340
rect 372724 316034 372752 336670
rect 372908 335354 372936 338014
rect 373000 338014 373060 338042
rect 373000 336734 373028 338014
rect 373322 337770 373350 338028
rect 373460 338014 373612 338042
rect 373736 338014 373888 338042
rect 374164 338014 374316 338042
rect 373322 337742 373396 337770
rect 372988 336728 373040 336734
rect 372988 336670 373040 336676
rect 372908 335326 373028 335354
rect 372896 326392 372948 326398
rect 372896 326334 372948 326340
rect 372804 326324 372856 326330
rect 372804 326266 372856 326272
rect 372632 316006 372752 316034
rect 372632 15910 372660 316006
rect 372712 313948 372764 313954
rect 372712 313890 372764 313896
rect 372724 16574 372752 313890
rect 372816 256018 372844 326266
rect 372908 286346 372936 326334
rect 373000 304298 373028 335326
rect 373368 330614 373396 337742
rect 373356 330608 373408 330614
rect 373356 330550 373408 330556
rect 373460 326398 373488 338014
rect 373448 326392 373500 326398
rect 373448 326334 373500 326340
rect 373736 326330 373764 338014
rect 374288 336326 374316 338014
rect 374380 338014 374440 338042
rect 374564 338014 374716 338042
rect 374840 338014 374992 338042
rect 375116 338014 375268 338042
rect 375484 338014 375544 338042
rect 375820 338014 375972 338042
rect 376096 338014 376248 338042
rect 374276 336320 374328 336326
rect 374276 336262 374328 336268
rect 374184 326392 374236 326398
rect 374184 326334 374236 326340
rect 373724 326324 373776 326330
rect 373724 326266 373776 326272
rect 374000 323604 374052 323610
rect 374000 323546 374052 323552
rect 372988 304292 373040 304298
rect 372988 304234 373040 304240
rect 372896 286340 372948 286346
rect 372896 286282 372948 286288
rect 372804 256012 372856 256018
rect 372804 255954 372856 255960
rect 372724 16546 372936 16574
rect 372620 15904 372672 15910
rect 372620 15846 372672 15852
rect 371884 4820 371936 4826
rect 371884 4762 371936 4768
rect 372908 480 372936 16546
rect 374012 3346 374040 323546
rect 374092 284980 374144 284986
rect 374092 284922 374144 284928
rect 374104 3466 374132 284922
rect 374196 254590 374224 326334
rect 374276 326324 374328 326330
rect 374276 326266 374328 326272
rect 374288 283626 374316 326266
rect 374380 284986 374408 338014
rect 374564 326398 374592 338014
rect 374552 326392 374604 326398
rect 374552 326334 374604 326340
rect 374840 323678 374868 338014
rect 375116 326330 375144 338014
rect 375380 326392 375432 326398
rect 375380 326334 375432 326340
rect 375104 326324 375156 326330
rect 375104 326266 375156 326272
rect 374828 323672 374880 323678
rect 374828 323614 374880 323620
rect 374368 284980 374420 284986
rect 374368 284922 374420 284928
rect 374276 283620 374328 283626
rect 374276 283562 374328 283568
rect 374184 254584 374236 254590
rect 374184 254526 374236 254532
rect 375392 253230 375420 326334
rect 375484 293282 375512 338014
rect 375944 329186 375972 338014
rect 376220 336734 376248 338014
rect 376312 338014 376372 338042
rect 376496 338014 376648 338042
rect 376924 338014 377076 338042
rect 376208 336728 376260 336734
rect 376208 336670 376260 336676
rect 375932 329180 375984 329186
rect 375932 329122 375984 329128
rect 376312 326398 376340 338014
rect 376496 327758 376524 338014
rect 377048 331226 377076 338014
rect 377140 338014 377200 338042
rect 377036 331220 377088 331226
rect 377036 331162 377088 331168
rect 377140 328250 377168 338014
rect 377462 337770 377490 338028
rect 377600 338014 377752 338042
rect 377876 338014 378028 338042
rect 378304 338014 378456 338042
rect 377462 337742 377536 337770
rect 377404 336728 377456 336734
rect 377404 336670 377456 336676
rect 377220 331220 377272 331226
rect 377220 331162 377272 331168
rect 376772 328222 377168 328250
rect 376484 327752 376536 327758
rect 376484 327694 376536 327700
rect 376300 326392 376352 326398
rect 376300 326334 376352 326340
rect 375472 293276 375524 293282
rect 375472 293218 375524 293224
rect 375380 253224 375432 253230
rect 375380 253166 375432 253172
rect 375380 25560 375432 25566
rect 375380 25502 375432 25508
rect 375392 16574 375420 25502
rect 376772 21418 376800 328222
rect 376944 326256 376996 326262
rect 376944 326198 376996 326204
rect 376852 326188 376904 326194
rect 376852 326130 376904 326136
rect 376864 251870 376892 326130
rect 376956 282198 376984 326198
rect 377232 324970 377260 331162
rect 377220 324964 377272 324970
rect 377220 324906 377272 324912
rect 377416 302938 377444 336670
rect 377508 336598 377536 337742
rect 377496 336592 377548 336598
rect 377496 336534 377548 336540
rect 377600 326262 377628 338014
rect 377588 326256 377640 326262
rect 377588 326198 377640 326204
rect 377876 326194 377904 338014
rect 378324 336728 378376 336734
rect 378324 336670 378376 336676
rect 378232 326392 378284 326398
rect 378232 326334 378284 326340
rect 378140 326324 378192 326330
rect 378140 326266 378192 326272
rect 377864 326188 377916 326194
rect 377864 326130 377916 326136
rect 377404 302932 377456 302938
rect 377404 302874 377456 302880
rect 376944 282192 376996 282198
rect 376944 282134 376996 282140
rect 376852 251864 376904 251870
rect 376852 251806 376904 251812
rect 376760 21412 376812 21418
rect 376760 21354 376812 21360
rect 375392 16546 376064 16574
rect 374092 3460 374144 3466
rect 374092 3402 374144 3408
rect 375288 3460 375340 3466
rect 375288 3402 375340 3408
rect 374012 3318 374132 3346
rect 374104 480 374132 3318
rect 375300 480 375328 3402
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 378152 14482 378180 326266
rect 378244 320958 378272 326334
rect 378232 320952 378284 320958
rect 378232 320894 378284 320900
rect 378232 307080 378284 307086
rect 378232 307022 378284 307028
rect 378244 16574 378272 307022
rect 378336 301510 378364 336670
rect 378428 335354 378456 338014
rect 378520 338014 378580 338042
rect 378704 338014 378856 338042
rect 378980 338014 379132 338042
rect 379256 338014 379408 338042
rect 379624 338014 379684 338042
rect 379808 338014 379960 338042
rect 380084 338014 380236 338042
rect 380360 338014 380512 338042
rect 378520 336734 378548 338014
rect 378508 336728 378560 336734
rect 378508 336670 378560 336676
rect 378704 335354 378732 338014
rect 378784 336388 378836 336394
rect 378784 336330 378836 336336
rect 378428 335326 378548 335354
rect 378520 322250 378548 335326
rect 378612 335326 378732 335354
rect 378508 322244 378560 322250
rect 378508 322186 378560 322192
rect 378612 321554 378640 335326
rect 378428 321526 378640 321554
rect 378428 305658 378456 321526
rect 378416 305652 378468 305658
rect 378416 305594 378468 305600
rect 378324 301504 378376 301510
rect 378324 301446 378376 301452
rect 378244 16546 378456 16574
rect 378140 14476 378192 14482
rect 378140 14418 378192 14424
rect 377680 4820 377732 4826
rect 377680 4762 377732 4768
rect 377692 480 377720 4762
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 378796 4554 378824 336330
rect 378980 326398 379008 338014
rect 378968 326392 379020 326398
rect 378968 326334 379020 326340
rect 379256 326330 379284 338014
rect 379520 326392 379572 326398
rect 379520 326334 379572 326340
rect 379244 326324 379296 326330
rect 379244 326266 379296 326272
rect 379532 250510 379560 326334
rect 379624 291854 379652 338014
rect 379808 326262 379836 338014
rect 379796 326256 379848 326262
rect 379796 326198 379848 326204
rect 380084 323610 380112 338014
rect 380360 326398 380388 338014
rect 380774 337770 380802 338028
rect 381064 338014 381216 338042
rect 380774 337742 380848 337770
rect 380820 334626 380848 337742
rect 380808 334620 380860 334626
rect 380808 334562 380860 334568
rect 380348 326392 380400 326398
rect 380348 326334 380400 326340
rect 381084 326392 381136 326398
rect 381084 326334 381136 326340
rect 380992 326324 381044 326330
rect 380992 326266 381044 326272
rect 380900 324148 380952 324154
rect 380900 324090 380952 324096
rect 380072 323604 380124 323610
rect 380072 323546 380124 323552
rect 379612 291848 379664 291854
rect 379612 291790 379664 291796
rect 379520 250504 379572 250510
rect 379520 250446 379572 250452
rect 380912 22778 380940 324090
rect 381004 249082 381032 326266
rect 381096 280838 381124 326334
rect 381188 300150 381216 338014
rect 381280 338014 381340 338042
rect 381464 338014 381616 338042
rect 381740 338014 381892 338042
rect 382016 338014 382168 338042
rect 382384 338014 382444 338042
rect 382568 338014 382720 338042
rect 382844 338014 382996 338042
rect 383120 338014 383272 338042
rect 383396 338014 383548 338042
rect 383764 338014 383824 338042
rect 384100 338014 384252 338042
rect 381280 324154 381308 338014
rect 381268 324148 381320 324154
rect 381268 324090 381320 324096
rect 381464 319462 381492 338014
rect 381740 326398 381768 338014
rect 381728 326392 381780 326398
rect 381728 326334 381780 326340
rect 382016 326330 382044 338014
rect 382384 336394 382412 338014
rect 382372 336388 382424 336394
rect 382372 336330 382424 336336
rect 382372 326528 382424 326534
rect 382372 326470 382424 326476
rect 382004 326324 382056 326330
rect 382004 326266 382056 326272
rect 382280 326324 382332 326330
rect 382280 326266 382332 326272
rect 381452 319456 381504 319462
rect 381452 319398 381504 319404
rect 381176 300144 381228 300150
rect 381176 300086 381228 300092
rect 381084 280832 381136 280838
rect 381084 280774 381136 280780
rect 380992 249076 381044 249082
rect 380992 249018 381044 249024
rect 382292 24138 382320 326266
rect 382384 47598 382412 326470
rect 382464 326392 382516 326398
rect 382464 326334 382516 326340
rect 382476 318102 382504 326334
rect 382464 318096 382516 318102
rect 382464 318038 382516 318044
rect 382568 279478 382596 338014
rect 382844 326330 382872 338014
rect 383120 326398 383148 338014
rect 383396 326534 383424 338014
rect 383384 326528 383436 326534
rect 383384 326470 383436 326476
rect 383108 326392 383160 326398
rect 383108 326334 383160 326340
rect 383660 326392 383712 326398
rect 383660 326334 383712 326340
rect 382832 326324 382884 326330
rect 382832 326266 382884 326272
rect 382464 279472 382516 279478
rect 382464 279414 382516 279420
rect 382556 279472 382608 279478
rect 382556 279414 382608 279420
rect 382372 47592 382424 47598
rect 382372 47534 382424 47540
rect 382280 24132 382332 24138
rect 382280 24074 382332 24080
rect 380900 22772 380952 22778
rect 380900 22714 380952 22720
rect 379520 15972 379572 15978
rect 379520 15914 379572 15920
rect 378784 4548 378836 4554
rect 378784 4490 378836 4496
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 379532 354 379560 15914
rect 381176 7608 381228 7614
rect 381176 7550 381228 7556
rect 381188 480 381216 7550
rect 382476 3602 382504 279414
rect 383672 247722 383700 326334
rect 383764 290494 383792 338014
rect 384224 331906 384252 338014
rect 384362 337770 384390 338028
rect 384500 338014 384652 338042
rect 384362 337742 384436 337770
rect 384212 331900 384264 331906
rect 384212 331842 384264 331848
rect 384408 329118 384436 337742
rect 384396 329112 384448 329118
rect 384396 329054 384448 329060
rect 384500 326398 384528 338014
rect 384914 337770 384942 338028
rect 385204 338014 385356 338042
rect 384914 337742 384988 337770
rect 384960 333266 384988 337742
rect 384948 333260 385000 333266
rect 384948 333202 385000 333208
rect 385328 326534 385356 338014
rect 385420 338014 385480 338042
rect 385604 338014 385756 338042
rect 385880 338014 386032 338042
rect 386156 338014 386308 338042
rect 386584 338014 386736 338042
rect 385316 326528 385368 326534
rect 385316 326470 385368 326476
rect 384488 326392 384540 326398
rect 384488 326334 384540 326340
rect 385040 326392 385092 326398
rect 385040 326334 385092 326340
rect 385052 298790 385080 326334
rect 385132 326324 385184 326330
rect 385132 326266 385184 326272
rect 385040 298784 385092 298790
rect 385040 298726 385092 298732
rect 383752 290488 383804 290494
rect 383752 290430 383804 290436
rect 385040 278044 385092 278050
rect 385040 277986 385092 277992
rect 383660 247716 383712 247722
rect 383660 247658 383712 247664
rect 382556 47728 382608 47734
rect 382556 47670 382608 47676
rect 382464 3596 382516 3602
rect 382464 3538 382516 3544
rect 382568 3482 382596 47670
rect 385052 16574 385080 277986
rect 385144 246362 385172 326266
rect 385420 323626 385448 338014
rect 385500 326528 385552 326534
rect 385500 326470 385552 326476
rect 385236 323598 385448 323626
rect 385236 269822 385264 323598
rect 385512 318794 385540 326470
rect 385328 318766 385540 318794
rect 385328 278050 385356 318766
rect 385604 316742 385632 338014
rect 385880 326398 385908 338014
rect 385868 326392 385920 326398
rect 385868 326334 385920 326340
rect 386156 326330 386184 338014
rect 386604 336728 386656 336734
rect 386604 336670 386656 336676
rect 386144 326324 386196 326330
rect 386144 326266 386196 326272
rect 386420 326324 386472 326330
rect 386420 326266 386472 326272
rect 385592 316736 385644 316742
rect 385592 316678 385644 316684
rect 385316 278044 385368 278050
rect 385316 277986 385368 277992
rect 385224 269816 385276 269822
rect 385224 269758 385276 269764
rect 385132 246356 385184 246362
rect 385132 246298 385184 246304
rect 385052 16546 386000 16574
rect 384764 4548 384816 4554
rect 384764 4490 384816 4496
rect 383568 3596 383620 3602
rect 383568 3538 383620 3544
rect 382384 3454 382596 3482
rect 382384 480 382412 3454
rect 383580 480 383608 3538
rect 384776 480 384804 4490
rect 385972 480 386000 16546
rect 386432 13122 386460 326266
rect 386512 324692 386564 324698
rect 386512 324634 386564 324640
rect 386524 182850 386552 324634
rect 386616 276690 386644 336670
rect 386708 335354 386736 338014
rect 386800 338014 386860 338042
rect 386984 338014 387136 338042
rect 387260 338014 387412 338042
rect 387536 338014 387688 338042
rect 387904 338014 387964 338042
rect 388180 338014 388240 338042
rect 388364 338014 388516 338042
rect 388640 338014 388792 338042
rect 388916 338014 389068 338042
rect 389192 338014 389344 338042
rect 389468 338014 389620 338042
rect 389744 338014 389896 338042
rect 390020 338014 390172 338042
rect 390296 338014 390448 338042
rect 390572 338014 390724 338042
rect 390848 338014 391000 338042
rect 391124 338014 391276 338042
rect 391400 338014 391552 338042
rect 391676 338014 391828 338042
rect 392044 338014 392104 338042
rect 392228 338014 392380 338042
rect 392504 338014 392656 338042
rect 392780 338014 392932 338042
rect 386800 336734 386828 338014
rect 386788 336728 386840 336734
rect 386788 336670 386840 336676
rect 386708 335326 386828 335354
rect 386696 326392 386748 326398
rect 386696 326334 386748 326340
rect 386708 313954 386736 326334
rect 386800 315314 386828 335326
rect 386984 326330 387012 338014
rect 387260 326398 387288 338014
rect 387248 326392 387300 326398
rect 387248 326334 387300 326340
rect 386972 326324 387024 326330
rect 386972 326266 387024 326272
rect 387536 324698 387564 338014
rect 387524 324692 387576 324698
rect 387524 324634 387576 324640
rect 387800 324352 387852 324358
rect 387800 324294 387852 324300
rect 386788 315308 386840 315314
rect 386788 315250 386840 315256
rect 386696 313948 386748 313954
rect 386696 313890 386748 313896
rect 386604 276684 386656 276690
rect 386604 276626 386656 276632
rect 386512 182844 386564 182850
rect 386512 182786 386564 182792
rect 386512 140072 386564 140078
rect 386512 140014 386564 140020
rect 386524 16574 386552 140014
rect 387812 17270 387840 324294
rect 387904 243574 387932 338014
rect 388076 326392 388128 326398
rect 388076 326334 388128 326340
rect 387984 323264 388036 323270
rect 387984 323206 388036 323212
rect 387996 275330 388024 323206
rect 388088 309806 388116 326334
rect 388180 311166 388208 338014
rect 388364 323270 388392 338014
rect 388640 324358 388668 338014
rect 388916 326398 388944 338014
rect 388904 326392 388956 326398
rect 388904 326334 388956 326340
rect 388628 324352 388680 324358
rect 388628 324294 388680 324300
rect 388352 323264 388404 323270
rect 388352 323206 388404 323212
rect 389192 320890 389220 338014
rect 389468 335354 389496 338014
rect 389376 335326 389496 335354
rect 389272 329452 389324 329458
rect 389272 329394 389324 329400
rect 389180 320884 389232 320890
rect 389180 320826 389232 320832
rect 389180 311296 389232 311302
rect 389180 311238 389232 311244
rect 388168 311160 388220 311166
rect 388168 311102 388220 311108
rect 388076 309800 388128 309806
rect 388076 309742 388128 309748
rect 387984 275324 388036 275330
rect 387984 275266 388036 275272
rect 387892 243568 387944 243574
rect 387892 243510 387944 243516
rect 387800 17264 387852 17270
rect 387800 17206 387852 17212
rect 389192 16574 389220 311238
rect 389284 90370 389312 329394
rect 389376 242214 389404 335326
rect 389456 330540 389508 330546
rect 389456 330482 389508 330488
rect 389468 273970 389496 330482
rect 389744 316034 389772 338014
rect 390020 330546 390048 338014
rect 390008 330540 390060 330546
rect 390008 330482 390060 330488
rect 390296 329458 390324 338014
rect 390572 330410 390600 338014
rect 390848 336682 390876 338014
rect 390664 336654 390876 336682
rect 390560 330404 390612 330410
rect 390560 330346 390612 330352
rect 390284 329452 390336 329458
rect 390284 329394 390336 329400
rect 390560 325100 390612 325106
rect 390560 325042 390612 325048
rect 389560 316006 389772 316034
rect 389560 308446 389588 316006
rect 389548 308440 389600 308446
rect 389548 308382 389600 308388
rect 389456 273964 389508 273970
rect 389456 273906 389508 273912
rect 389364 242208 389416 242214
rect 389364 242150 389416 242156
rect 389272 90364 389324 90370
rect 389272 90306 389324 90312
rect 386524 16546 386736 16574
rect 389192 16546 389496 16574
rect 386420 13116 386472 13122
rect 386420 13058 386472 13064
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 378846 -960 378958 326
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 386708 354 386736 16546
rect 387800 13184 387852 13190
rect 387800 13126 387852 13132
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 13126
rect 389468 480 389496 16546
rect 390572 3466 390600 325042
rect 390664 297430 390692 336654
rect 391124 335354 391152 338014
rect 390756 335326 391152 335354
rect 390652 297424 390704 297430
rect 390652 297366 390704 297372
rect 390652 271176 390704 271182
rect 390652 271118 390704 271124
rect 390560 3460 390612 3466
rect 390560 3402 390612 3408
rect 390664 480 390692 271118
rect 390756 171834 390784 335326
rect 390836 330540 390888 330546
rect 390836 330482 390888 330488
rect 390848 271182 390876 330482
rect 391400 316034 391428 338014
rect 391676 330546 391704 338014
rect 392044 335442 392072 338014
rect 392032 335436 392084 335442
rect 392032 335378 392084 335384
rect 391664 330540 391716 330546
rect 391664 330482 391716 330488
rect 391940 330540 391992 330546
rect 391940 330482 391992 330488
rect 390940 316006 391428 316034
rect 390940 307086 390968 316006
rect 390928 307080 390980 307086
rect 390928 307022 390980 307028
rect 390836 271176 390888 271182
rect 390836 271118 390888 271124
rect 390744 171828 390796 171834
rect 390744 171770 390796 171776
rect 391952 3466 391980 330482
rect 392032 330472 392084 330478
rect 392032 330414 392084 330420
rect 391848 3460 391900 3466
rect 391848 3402 391900 3408
rect 391940 3460 391992 3466
rect 391940 3402 391992 3408
rect 391860 480 391888 3402
rect 392044 3369 392072 330414
rect 392228 316034 392256 338014
rect 392504 330546 392532 338014
rect 392492 330540 392544 330546
rect 392492 330482 392544 330488
rect 392780 330478 392808 338014
rect 400862 337991 400918 338000
rect 399484 336592 399536 336598
rect 399484 336534 399536 336540
rect 395344 336524 395396 336530
rect 395344 336466 395396 336472
rect 393964 335436 394016 335442
rect 393964 335378 394016 335384
rect 392768 330472 392820 330478
rect 392768 330414 392820 330420
rect 392136 316006 392256 316034
rect 392136 3602 392164 316006
rect 393976 240786 394004 335378
rect 394700 322380 394752 322386
rect 394700 322322 394752 322328
rect 393964 240780 394016 240786
rect 393964 240722 394016 240728
rect 393320 26920 393372 26926
rect 393320 26862 393372 26868
rect 393332 16574 393360 26862
rect 393332 16546 394280 16574
rect 393044 8968 393096 8974
rect 393044 8910 393096 8916
rect 392124 3596 392176 3602
rect 392124 3538 392176 3544
rect 392030 3360 392086 3369
rect 392030 3295 392086 3304
rect 393056 480 393084 8910
rect 394252 480 394280 16546
rect 394712 6914 394740 322322
rect 395356 7614 395384 336466
rect 396724 336456 396776 336462
rect 396724 336398 396776 336404
rect 395434 334656 395490 334665
rect 395434 334591 395490 334600
rect 395448 233238 395476 334591
rect 396080 332036 396132 332042
rect 396080 331978 396132 331984
rect 395436 233232 395488 233238
rect 395436 233174 395488 233180
rect 395344 7608 395396 7614
rect 395344 7550 395396 7556
rect 394712 6886 395384 6914
rect 395356 480 395384 6886
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 331978
rect 396736 4826 396764 336398
rect 396814 333296 396870 333305
rect 396814 333231 396870 333240
rect 396828 325650 396856 333231
rect 396816 325644 396868 325650
rect 396816 325586 396868 325592
rect 398840 316872 398892 316878
rect 398840 316814 398892 316820
rect 397460 28280 397512 28286
rect 397460 28222 397512 28228
rect 397472 16574 397500 28222
rect 397472 16546 397776 16574
rect 396724 4820 396776 4826
rect 396724 4762 396776 4768
rect 397748 480 397776 16546
rect 398852 3074 398880 316814
rect 398932 17332 398984 17338
rect 398932 17274 398984 17280
rect 398944 3194 398972 17274
rect 399496 10334 399524 336534
rect 400220 86284 400272 86290
rect 400220 86226 400272 86232
rect 400232 16574 400260 86226
rect 400876 85542 400904 337991
rect 407764 336388 407816 336394
rect 407764 336330 407816 336336
rect 407120 330676 407172 330682
rect 407120 330618 407172 330624
rect 405002 327720 405058 327729
rect 405002 327655 405058 327664
rect 401600 321020 401652 321026
rect 401600 320962 401652 320968
rect 400864 85536 400916 85542
rect 400864 85478 400916 85484
rect 401612 16574 401640 320962
rect 402980 309936 403032 309942
rect 402980 309878 403032 309884
rect 402992 16574 403020 309878
rect 405016 179382 405044 327655
rect 405740 319592 405792 319598
rect 405740 319534 405792 319540
rect 405004 179376 405056 179382
rect 405004 179318 405056 179324
rect 404360 178696 404412 178702
rect 404360 178638 404412 178644
rect 400232 16546 400904 16574
rect 401612 16546 402560 16574
rect 402992 16546 403664 16574
rect 399484 10328 399536 10334
rect 399484 10270 399536 10276
rect 398932 3188 398984 3194
rect 398932 3130 398984 3136
rect 400128 3188 400180 3194
rect 400128 3130 400180 3136
rect 398852 3046 398972 3074
rect 398944 480 398972 3046
rect 400140 480 400168 3130
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 16546
rect 402532 480 402560 16546
rect 403636 480 403664 16546
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 178638
rect 405752 16574 405780 319534
rect 405752 16546 406056 16574
rect 406028 480 406056 16546
rect 407132 3074 407160 330618
rect 407212 29640 407264 29646
rect 407212 29582 407264 29588
rect 407224 3194 407252 29582
rect 407776 11762 407804 336330
rect 410524 336320 410576 336326
rect 410524 336262 410576 336268
rect 407854 326360 407910 326369
rect 407854 326295 407910 326304
rect 407868 259418 407896 326295
rect 408500 325032 408552 325038
rect 408500 324974 408552 324980
rect 407856 259412 407908 259418
rect 407856 259354 407908 259360
rect 408512 16574 408540 324974
rect 409880 308508 409932 308514
rect 409880 308450 409932 308456
rect 408512 16546 409184 16574
rect 407764 11756 407816 11762
rect 407764 11698 407816 11704
rect 407212 3188 407264 3194
rect 407212 3130 407264 3136
rect 408408 3188 408460 3194
rect 408408 3130 408460 3136
rect 407132 3046 407252 3074
rect 407224 480 407252 3046
rect 408420 480 408448 3130
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 409892 6914 409920 308450
rect 410536 8974 410564 336262
rect 412640 323740 412692 323746
rect 412640 323682 412692 323688
rect 411904 11824 411956 11830
rect 411904 11766 411956 11772
rect 410524 8968 410576 8974
rect 410524 8910 410576 8916
rect 409892 6886 410840 6914
rect 410812 480 410840 6886
rect 411916 480 411944 11766
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 323682
rect 413388 20670 413416 451246
rect 414020 272536 414072 272542
rect 414020 272478 414072 272484
rect 413376 20664 413428 20670
rect 413376 20606 413428 20612
rect 414032 16574 414060 272478
rect 414124 137290 414152 457438
rect 414112 137284 414164 137290
rect 414112 137226 414164 137232
rect 414676 86970 414704 458390
rect 416056 353258 416084 458730
rect 416044 353252 416096 353258
rect 416044 353194 416096 353200
rect 416780 312588 416832 312594
rect 416780 312530 416832 312536
rect 415400 305788 415452 305794
rect 415400 305730 415452 305736
rect 414664 86964 414716 86970
rect 414664 86906 414716 86912
rect 414032 16546 414336 16574
rect 414308 480 414336 16546
rect 415412 3262 415440 305730
rect 416792 16574 416820 312530
rect 417436 126954 417464 461246
rect 418804 458584 418856 458590
rect 418804 458526 418856 458532
rect 418160 258732 418212 258738
rect 418160 258674 418212 258680
rect 417424 126948 417476 126954
rect 417424 126890 417476 126896
rect 418172 16574 418200 258674
rect 418816 167006 418844 458526
rect 419540 318232 419592 318238
rect 419540 318174 419592 318180
rect 418804 167000 418856 167006
rect 418804 166942 418856 166948
rect 419552 16574 419580 318174
rect 420920 269884 420972 269890
rect 420920 269826 420972 269832
rect 416792 16546 417464 16574
rect 418172 16546 418568 16574
rect 419552 16546 420224 16574
rect 415492 4888 415544 4894
rect 415492 4830 415544 4836
rect 415400 3256 415452 3262
rect 415400 3198 415452 3204
rect 415504 480 415532 4830
rect 416688 3256 416740 3262
rect 416688 3198 416740 3204
rect 416700 480 416728 3198
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 420196 480 420224 16546
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 269826
rect 421576 206990 421604 462606
rect 422956 245614 422984 462742
rect 427084 462528 427136 462534
rect 427084 462470 427136 462476
rect 424324 462460 424376 462466
rect 424324 462402 424376 462408
rect 423680 316804 423732 316810
rect 423680 316746 423732 316752
rect 422944 245608 422996 245614
rect 422944 245550 422996 245556
rect 422300 244928 422352 244934
rect 422300 244870 422352 244876
rect 421564 206984 421616 206990
rect 421564 206926 421616 206932
rect 422312 16574 422340 244870
rect 422312 16546 422616 16574
rect 422588 480 422616 16546
rect 423692 3330 423720 316746
rect 423772 304360 423824 304366
rect 423772 304302 423824 304308
rect 423680 3324 423732 3330
rect 423680 3266 423732 3272
rect 423784 480 423812 304302
rect 424336 73166 424364 462402
rect 426440 329248 426492 329254
rect 426440 329190 426492 329196
rect 424324 73160 424376 73166
rect 424324 73102 424376 73108
rect 426452 16574 426480 329190
rect 427096 113150 427124 462470
rect 428464 461236 428516 461242
rect 428464 461178 428516 461184
rect 427820 307148 427872 307154
rect 427820 307090 427872 307096
rect 427084 113144 427136 113150
rect 427084 113086 427136 113092
rect 427832 16574 427860 307090
rect 428476 193186 428504 461178
rect 431224 458516 431276 458522
rect 431224 458458 431276 458464
rect 430580 315444 430632 315450
rect 430580 315386 430632 315392
rect 428464 193180 428516 193186
rect 428464 193122 428516 193128
rect 430592 16574 430620 315386
rect 431236 273222 431264 458458
rect 432604 456884 432656 456890
rect 432604 456826 432656 456832
rect 432616 379506 432644 456826
rect 432604 379500 432656 379506
rect 432604 379442 432656 379448
rect 435376 365702 435404 464034
rect 457444 463820 457496 463826
rect 457444 463762 457496 463768
rect 454684 462596 454736 462602
rect 454684 462538 454736 462544
rect 454696 405686 454724 462538
rect 457456 431934 457484 463762
rect 462332 460834 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 462320 460828 462372 460834
rect 462320 460770 462372 460776
rect 477512 460766 477540 702406
rect 494072 472666 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 494060 472660 494112 472666
rect 494060 472602 494112 472608
rect 477500 460760 477552 460766
rect 477500 460702 477552 460708
rect 527192 460630 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 527180 460624 527232 460630
rect 527180 460566 527232 460572
rect 542372 460562 542400 702406
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670812 580224 670818
rect 580172 670754 580224 670760
rect 580184 670721 580212 670754
rect 580170 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 567936 461032 567988 461038
rect 567936 460974 567988 460980
rect 542360 460556 542412 460562
rect 542360 460498 542412 460504
rect 457444 431928 457496 431934
rect 457444 431870 457496 431876
rect 454684 405680 454736 405686
rect 454684 405622 454736 405628
rect 435364 365696 435416 365702
rect 435364 365638 435416 365644
rect 432602 337512 432658 337521
rect 432602 337447 432658 337456
rect 432052 319524 432104 319530
rect 432052 319466 432104 319472
rect 431224 273216 431276 273222
rect 431224 273158 431276 273164
rect 426452 16546 426848 16574
rect 427832 16546 428504 16574
rect 430592 16546 430896 16574
rect 424968 3324 425020 3330
rect 424968 3266 425020 3272
rect 424980 480 425008 3266
rect 426164 3120 426216 3126
rect 426164 3062 426216 3068
rect 426176 480 426204 3062
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 426820 354 426848 16546
rect 428476 480 428504 16546
rect 429660 3188 429712 3194
rect 429660 3130 429712 3136
rect 429672 480 429700 3130
rect 430868 480 430896 16546
rect 432064 480 432092 319466
rect 432616 219434 432644 337447
rect 436100 336252 436152 336258
rect 436100 336194 436152 336200
rect 434720 311228 434772 311234
rect 434720 311170 434772 311176
rect 433340 303000 433392 303006
rect 433340 302942 433392 302948
rect 432604 219428 432656 219434
rect 432604 219370 432656 219376
rect 433352 16574 433380 302942
rect 434732 16574 434760 311170
rect 436112 16574 436140 336194
rect 443000 336184 443052 336190
rect 443000 336126 443052 336132
rect 438860 334756 438912 334762
rect 438860 334698 438912 334704
rect 437480 301572 437532 301578
rect 437480 301514 437532 301520
rect 433352 16546 434024 16574
rect 434732 16546 435128 16574
rect 436112 16546 436784 16574
rect 433248 3392 433300 3398
rect 433248 3334 433300 3340
rect 433260 480 433288 3334
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 16546
rect 436756 480 436784 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 301514
rect 438872 16574 438900 334698
rect 441620 333396 441672 333402
rect 441620 333338 441672 333344
rect 440332 300212 440384 300218
rect 440332 300154 440384 300160
rect 438872 16546 439176 16574
rect 439148 480 439176 16546
rect 440240 4140 440292 4146
rect 440240 4082 440292 4088
rect 440252 2122 440280 4082
rect 440344 3398 440372 300154
rect 441632 16574 441660 333338
rect 443012 16574 443040 336126
rect 449900 336116 449952 336122
rect 449900 336058 449952 336064
rect 448520 327820 448572 327826
rect 448520 327762 448572 327768
rect 444380 298852 444432 298858
rect 444380 298794 444432 298800
rect 444392 16574 444420 298794
rect 445760 268388 445812 268394
rect 445760 268330 445812 268336
rect 441632 16546 442672 16574
rect 443012 16546 443408 16574
rect 444392 16546 445064 16574
rect 440332 3392 440384 3398
rect 440332 3334 440384 3340
rect 441528 3392 441580 3398
rect 441528 3334 441580 3340
rect 440252 2094 440372 2122
rect 440344 480 440372 2094
rect 441540 480 441568 3334
rect 442644 480 442672 16546
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 16546
rect 445036 480 445064 16546
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 445772 354 445800 268330
rect 447416 4072 447468 4078
rect 447416 4014 447468 4020
rect 447428 480 447456 4014
rect 448532 3210 448560 327762
rect 448612 318164 448664 318170
rect 448612 318106 448664 318112
rect 448624 3398 448652 318106
rect 449912 16574 449940 336058
rect 456800 336048 456852 336054
rect 456800 335990 456852 335996
rect 451280 297492 451332 297498
rect 451280 297434 451332 297440
rect 451292 16574 451320 297434
rect 455420 296064 455472 296070
rect 455420 296006 455472 296012
rect 452660 267028 452712 267034
rect 452660 266970 452712 266976
rect 452672 16574 452700 266970
rect 455432 16574 455460 296006
rect 449912 16546 450952 16574
rect 451292 16546 451688 16574
rect 452672 16546 453344 16574
rect 455432 16546 455736 16574
rect 448612 3392 448664 3398
rect 448612 3334 448664 3340
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 448532 3182 448652 3210
rect 448624 480 448652 3182
rect 449820 480 449848 3334
rect 450924 480 450952 16546
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 453316 480 453344 16546
rect 454500 4004 454552 4010
rect 454500 3946 454552 3952
rect 454512 480 454540 3946
rect 455708 480 455736 16546
rect 456812 1698 456840 335990
rect 480260 334688 480312 334694
rect 480260 334630 480312 334636
rect 462320 326460 462372 326466
rect 462320 326402 462372 326408
rect 459560 309868 459612 309874
rect 459560 309810 459612 309816
rect 458180 294704 458232 294710
rect 458180 294646 458232 294652
rect 456892 265668 456944 265674
rect 456892 265610 456944 265616
rect 456800 1692 456852 1698
rect 456800 1634 456852 1640
rect 456904 480 456932 265610
rect 458192 16574 458220 294646
rect 459572 16574 459600 309810
rect 458192 16546 459232 16574
rect 459572 16546 459968 16574
rect 458088 1692 458140 1698
rect 458088 1634 458140 1640
rect 458100 480 458128 1634
rect 459204 480 459232 16546
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 461584 3936 461636 3942
rect 461584 3878 461636 3884
rect 461596 480 461624 3878
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 326402
rect 469220 322312 469272 322318
rect 469220 322254 469272 322260
rect 466460 315376 466512 315382
rect 466460 315318 466512 315324
rect 465172 293344 465224 293350
rect 465172 293286 465224 293292
rect 463700 264240 463752 264246
rect 463700 264182 463752 264188
rect 463712 16574 463740 264182
rect 465184 16574 465212 293286
rect 466472 16574 466500 315318
rect 469232 16574 469260 322254
rect 473360 305720 473412 305726
rect 473360 305662 473412 305668
rect 470600 295996 470652 296002
rect 470600 295938 470652 295944
rect 463712 16546 464016 16574
rect 465184 16546 465856 16574
rect 466472 16546 467512 16574
rect 469232 16546 469904 16574
rect 463988 480 464016 16546
rect 465172 3868 465224 3874
rect 465172 3810 465224 3816
rect 465184 480 465212 3810
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 354 465856 16546
rect 467484 480 467512 16546
rect 468668 3800 468720 3806
rect 468668 3742 468720 3748
rect 468680 480 468708 3742
rect 469876 480 469904 16546
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 354 470640 295938
rect 473372 6914 473400 305662
rect 476120 291916 476172 291922
rect 476120 291858 476172 291864
rect 473452 262880 473504 262886
rect 473452 262822 473504 262828
rect 473464 16574 473492 262822
rect 476132 16574 476160 291858
rect 477500 261520 477552 261526
rect 477500 261462 477552 261468
rect 477512 16574 477540 261462
rect 480272 16574 480300 334630
rect 529940 334620 529992 334626
rect 529940 334562 529992 334568
rect 494060 333328 494112 333334
rect 494060 333270 494112 333276
rect 489920 331968 489972 331974
rect 489920 331910 489972 331916
rect 481640 314016 481692 314022
rect 481640 313958 481692 313964
rect 473464 16546 474136 16574
rect 476132 16546 476528 16574
rect 477512 16546 478184 16574
rect 480272 16546 480576 16574
rect 473372 6886 473492 6914
rect 472256 3732 472308 3738
rect 472256 3674 472308 3680
rect 472268 480 472296 3674
rect 473464 480 473492 6886
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 16546
rect 475752 3664 475804 3670
rect 475752 3606 475804 3612
rect 475764 480 475792 3606
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 478156 480 478184 16546
rect 479340 3528 479392 3534
rect 479340 3470 479392 3476
rect 479352 480 479380 3470
rect 480548 480 480576 16546
rect 481652 6914 481680 313958
rect 484400 290556 484452 290562
rect 484400 290498 484452 290504
rect 481732 18624 481784 18630
rect 481732 18566 481784 18572
rect 481744 16574 481772 18566
rect 484412 16574 484440 290498
rect 488540 289128 488592 289134
rect 488540 289070 488592 289076
rect 485780 260160 485832 260166
rect 485780 260102 485832 260108
rect 485792 16574 485820 260102
rect 488552 16574 488580 289070
rect 481744 16546 482416 16574
rect 484412 16546 484808 16574
rect 485792 16546 486464 16574
rect 488552 16546 488856 16574
rect 481652 6886 481772 6914
rect 481744 480 481772 6886
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 354 482416 16546
rect 484032 4820 484084 4826
rect 484032 4762 484084 4768
rect 484044 480 484072 4762
rect 482806 354 482918 480
rect 482388 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 486436 480 486464 16546
rect 487620 7608 487672 7614
rect 487620 7550 487672 7556
rect 487632 480 487660 7550
rect 488828 480 488856 16546
rect 489932 3534 489960 331910
rect 490012 294636 490064 294642
rect 490012 294578 490064 294584
rect 489920 3528 489972 3534
rect 489920 3470 489972 3476
rect 490024 3346 490052 294578
rect 491300 287700 491352 287706
rect 491300 287642 491352 287648
rect 491312 16574 491340 287642
rect 492680 257372 492732 257378
rect 492680 257314 492732 257320
rect 492692 16574 492720 257314
rect 494072 16574 494100 333270
rect 498200 330608 498252 330614
rect 498200 330550 498252 330556
rect 495440 304292 495492 304298
rect 495440 304234 495492 304240
rect 491312 16546 492352 16574
rect 492692 16546 493088 16574
rect 494072 16546 494744 16574
rect 490748 3528 490800 3534
rect 490748 3470 490800 3476
rect 489932 3318 490052 3346
rect 489932 480 489960 3318
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490760 354 490788 3470
rect 492324 480 492352 16546
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494716 480 494744 16546
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 304234
rect 497096 15904 497148 15910
rect 497096 15846 497148 15852
rect 497108 480 497136 15846
rect 498212 480 498240 330550
rect 507860 329180 507912 329186
rect 507860 329122 507912 329128
rect 505100 323672 505152 323678
rect 505100 323614 505152 323620
rect 498292 286340 498344 286346
rect 498292 286282 498344 286288
rect 498304 16574 498332 286282
rect 502340 284980 502392 284986
rect 502340 284922 502392 284928
rect 499580 256012 499632 256018
rect 499580 255954 499632 255960
rect 499592 16574 499620 255954
rect 502352 16574 502380 284922
rect 503720 254584 503772 254590
rect 503720 254526 503772 254532
rect 498304 16546 498976 16574
rect 499592 16546 500632 16574
rect 502352 16546 503024 16574
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 354 498976 16546
rect 500604 480 500632 16546
rect 501788 8968 501840 8974
rect 501788 8910 501840 8916
rect 501800 480 501828 8910
rect 502996 480 503024 16546
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 354 503760 254526
rect 505112 16574 505140 323614
rect 506480 293276 506532 293282
rect 506480 293218 506532 293224
rect 505112 16546 505416 16574
rect 505388 480 505416 16546
rect 506492 3534 506520 293218
rect 506572 283620 506624 283626
rect 506572 283562 506624 283568
rect 506480 3528 506532 3534
rect 506480 3470 506532 3476
rect 506584 3346 506612 283562
rect 507872 16574 507900 329122
rect 512000 327752 512052 327758
rect 512000 327694 512052 327700
rect 509240 302932 509292 302938
rect 509240 302874 509292 302880
rect 509252 16574 509280 302874
rect 510620 253224 510672 253230
rect 510620 253166 510672 253172
rect 510632 16574 510660 253166
rect 507872 16546 508912 16574
rect 509252 16546 509648 16574
rect 510632 16546 511304 16574
rect 507308 3528 507360 3534
rect 507308 3470 507360 3476
rect 506492 3318 506612 3346
rect 506492 480 506520 3318
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507320 354 507348 3470
rect 508884 480 508912 16546
rect 507646 354 507758 480
rect 507320 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 511276 480 511304 16546
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 327694
rect 525800 326392 525852 326398
rect 525800 326334 525852 326340
rect 513380 324964 513432 324970
rect 513380 324906 513432 324912
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 324906
rect 518900 322244 518952 322250
rect 518900 322186 518952 322192
rect 516140 282192 516192 282198
rect 516140 282134 516192 282140
rect 514760 21412 514812 21418
rect 514760 21354 514812 21360
rect 514772 480 514800 21354
rect 516152 16574 516180 282134
rect 517520 251864 517572 251870
rect 517520 251806 517572 251812
rect 517532 16574 517560 251806
rect 518912 16574 518940 322186
rect 523040 320952 523092 320958
rect 523040 320894 523092 320900
rect 521660 305652 521712 305658
rect 521660 305594 521712 305600
rect 520280 301504 520332 301510
rect 520280 301446 520332 301452
rect 516152 16546 517192 16574
rect 517532 16546 517928 16574
rect 518912 16546 519584 16574
rect 515496 10328 515548 10334
rect 515496 10270 515548 10276
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515508 354 515536 10270
rect 517164 480 517192 16546
rect 515926 354 516038 480
rect 515508 326 516038 354
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519556 480 519584 16546
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 301446
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 305594
rect 523052 480 523080 320894
rect 524420 291848 524472 291854
rect 524420 291790 524472 291796
rect 524432 16574 524460 291790
rect 525812 16574 525840 326334
rect 527180 323604 527232 323610
rect 527180 323546 527232 323552
rect 527192 16574 527220 323546
rect 528560 250504 528612 250510
rect 528560 250446 528612 250452
rect 524432 16546 525472 16574
rect 525812 16546 526208 16574
rect 527192 16546 527864 16574
rect 523776 14476 523828 14482
rect 523776 14418 523828 14424
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523788 354 523816 14418
rect 525444 480 525472 16546
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527836 480 527864 16546
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 250446
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 334562
rect 547880 333260 547932 333266
rect 547880 333202 547932 333208
rect 543740 331900 543792 331906
rect 543740 331842 543792 331848
rect 532700 319456 532752 319462
rect 532700 319398 532752 319404
rect 531320 300144 531372 300150
rect 531320 300086 531372 300092
rect 531332 480 531360 300086
rect 531412 22772 531464 22778
rect 531412 22714 531464 22720
rect 531424 16574 531452 22714
rect 532712 16574 532740 319398
rect 539600 318096 539652 318102
rect 539600 318038 539652 318044
rect 534080 280832 534132 280838
rect 534080 280774 534132 280780
rect 534092 16574 534120 280774
rect 538220 279472 538272 279478
rect 538220 279414 538272 279420
rect 535460 249076 535512 249082
rect 535460 249018 535512 249024
rect 535472 16574 535500 249018
rect 531424 16546 532096 16574
rect 532712 16546 533752 16574
rect 534092 16546 534488 16574
rect 535472 16546 536144 16574
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532068 354 532096 16546
rect 533724 480 533752 16546
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536116 480 536144 16546
rect 537208 11756 537260 11762
rect 537208 11698 537260 11704
rect 537220 480 537248 11698
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 279414
rect 539612 3534 539640 318038
rect 542360 290488 542412 290494
rect 542360 290430 542412 290436
rect 540980 47592 541032 47598
rect 540980 47534 541032 47540
rect 539692 24132 539744 24138
rect 539692 24074 539744 24080
rect 539600 3528 539652 3534
rect 539600 3470 539652 3476
rect 539704 3346 539732 24074
rect 540992 16574 541020 47534
rect 542372 16574 542400 290430
rect 543752 16574 543780 331842
rect 545120 329112 545172 329118
rect 545120 329054 545172 329060
rect 545132 16574 545160 329054
rect 546500 247716 546552 247722
rect 546500 247658 546552 247664
rect 540992 16546 542032 16574
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 545132 16546 545528 16574
rect 540428 3528 540480 3534
rect 540428 3470 540480 3476
rect 539612 3318 539732 3346
rect 539612 480 539640 3318
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540440 354 540468 3470
rect 542004 480 542032 16546
rect 540766 354 540878 480
rect 540440 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545500 480 545528 16546
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 247658
rect 547892 480 547920 333202
rect 565820 320884 565872 320890
rect 565820 320826 565872 320832
rect 550640 316736 550692 316742
rect 550640 316678 550692 316684
rect 547972 278044 548024 278050
rect 547972 277986 548024 277992
rect 547984 16574 548012 277986
rect 549260 269816 549312 269822
rect 549260 269758 549312 269764
rect 549272 16574 549300 269758
rect 550652 16574 550680 316678
rect 554780 315308 554832 315314
rect 554780 315250 554832 315256
rect 552020 298784 552072 298790
rect 552020 298726 552072 298732
rect 552032 16574 552060 298726
rect 553400 246356 553452 246362
rect 553400 246298 553452 246304
rect 553412 16574 553440 246298
rect 554042 164928 554098 164937
rect 554042 164863 554098 164872
rect 554056 153202 554084 164863
rect 554044 153196 554096 153202
rect 554044 153138 554096 153144
rect 547984 16546 548656 16574
rect 549272 16546 550312 16574
rect 550652 16546 551048 16574
rect 552032 16546 552704 16574
rect 553412 16546 553808 16574
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548628 354 548656 16546
rect 550284 480 550312 16546
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 552676 480 552704 16546
rect 553780 480 553808 16546
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 315250
rect 557540 313948 557592 313954
rect 557540 313890 557592 313896
rect 556160 276684 556212 276690
rect 556160 276626 556212 276632
rect 556172 480 556200 276626
rect 557552 16574 557580 313890
rect 561680 311160 561732 311166
rect 561680 311102 561732 311108
rect 560300 243568 560352 243574
rect 560300 243510 560352 243516
rect 558920 182844 558972 182850
rect 558920 182786 558972 182792
rect 558932 16574 558960 182786
rect 560312 16574 560340 243510
rect 561692 16574 561720 311102
rect 564440 309800 564492 309806
rect 564440 309742 564492 309748
rect 563060 275324 563112 275330
rect 563060 275266 563112 275272
rect 557552 16546 558592 16574
rect 558932 16546 559328 16574
rect 560312 16546 560432 16574
rect 561692 16546 562088 16574
rect 556896 13116 556948 13122
rect 556896 13058 556948 13064
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 556908 354 556936 13058
rect 558564 480 558592 16546
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 562060 480 562088 16546
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 275266
rect 564452 3534 564480 309742
rect 564532 17264 564584 17270
rect 564532 17206 564584 17212
rect 564440 3528 564492 3534
rect 564440 3470 564492 3476
rect 564544 3346 564572 17206
rect 565832 16574 565860 320826
rect 567844 308440 567896 308446
rect 567844 308382 567896 308388
rect 567200 242208 567252 242214
rect 567200 242150 567252 242156
rect 567212 16574 567240 242150
rect 565832 16546 566872 16574
rect 567212 16546 567608 16574
rect 565268 3528 565320 3534
rect 565268 3470 565320 3476
rect 564452 3318 564572 3346
rect 564452 480 564480 3318
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565280 354 565308 3470
rect 566844 480 566872 16546
rect 565606 354 565718 480
rect 565280 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 567856 3534 567884 308382
rect 567948 299470 567976 460974
rect 580356 458856 580408 458862
rect 580356 458798 580408 458804
rect 580264 458312 580316 458318
rect 580264 458254 580316 458260
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 579620 431928 579672 431934
rect 579620 431870 579672 431876
rect 579632 431633 579660 431870
rect 579618 431624 579674 431633
rect 579618 431559 579674 431568
rect 579620 405680 579672 405686
rect 579620 405622 579672 405628
rect 579632 404977 579660 405622
rect 579618 404968 579674 404977
rect 579618 404903 579674 404912
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 571984 330540 572036 330546
rect 571984 330482 572036 330488
rect 567936 299464 567988 299470
rect 567936 299406 567988 299412
rect 569960 273964 570012 273970
rect 569960 273906 570012 273912
rect 569972 16574 570000 273906
rect 570604 90364 570656 90370
rect 570604 90306 570656 90312
rect 569972 16546 570368 16574
rect 567844 3528 567896 3534
rect 567844 3470 567896 3476
rect 569132 3528 569184 3534
rect 569132 3470 569184 3476
rect 569144 480 569172 3470
rect 570340 480 570368 16546
rect 570616 3534 570644 90306
rect 571996 3534 572024 330482
rect 579896 325644 579948 325650
rect 579896 325586 579948 325592
rect 579908 325281 579936 325586
rect 579894 325272 579950 325281
rect 579894 325207 579950 325216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 575480 307080 575532 307086
rect 575480 307022 575532 307028
rect 572076 297424 572128 297430
rect 572076 297366 572128 297372
rect 570604 3528 570656 3534
rect 570604 3470 570656 3476
rect 571524 3528 571576 3534
rect 571524 3470 571576 3476
rect 571984 3528 572036 3534
rect 571984 3470 572036 3476
rect 571536 480 571564 3470
rect 572088 3398 572116 297366
rect 574744 271176 574796 271182
rect 574744 271118 574796 271124
rect 574100 171828 574152 171834
rect 574100 171770 574152 171776
rect 574112 16574 574140 171770
rect 574112 16546 574692 16574
rect 572720 3528 572772 3534
rect 572720 3470 572772 3476
rect 574664 3482 574692 16546
rect 574756 3874 574784 271118
rect 575492 16574 575520 307022
rect 579620 299464 579672 299470
rect 579620 299406 579672 299412
rect 579632 298761 579660 299406
rect 579618 298752 579674 298761
rect 579618 298687 579674 298696
rect 579896 273216 579948 273222
rect 579896 273158 579948 273164
rect 579908 272241 579936 273158
rect 579894 272232 579950 272241
rect 579894 272167 579950 272176
rect 579804 259412 579856 259418
rect 579804 259354 579856 259360
rect 579816 258913 579844 259354
rect 579802 258904 579858 258913
rect 579802 258839 579858 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 578240 240780 578292 240786
rect 578240 240722 578292 240728
rect 578252 16574 578280 240722
rect 580172 233232 580224 233238
rect 580172 233174 580224 233180
rect 580184 232393 580212 233174
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 579896 219428 579948 219434
rect 579896 219370 579948 219376
rect 579908 219065 579936 219370
rect 579894 219056 579950 219065
rect 579894 218991 579950 219000
rect 580172 206984 580224 206990
rect 580172 206926 580224 206932
rect 580184 205737 580212 206926
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 579988 179376 580040 179382
rect 579988 179318 580040 179324
rect 580000 179217 580028 179318
rect 579986 179208 580042 179217
rect 579986 179143 580042 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 579804 153196 579856 153202
rect 579804 153138 579856 153144
rect 579816 152697 579844 153138
rect 579802 152688 579858 152697
rect 579802 152623 579858 152632
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 580172 113144 580224 113150
rect 580172 113086 580224 113092
rect 580184 112849 580212 113086
rect 580170 112840 580226 112849
rect 580170 112775 580226 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 579988 73160 580040 73166
rect 579988 73102 580040 73108
rect 580000 73001 580028 73102
rect 579986 72992 580042 73001
rect 579986 72927 580042 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580276 46345 580304 458254
rect 580368 418305 580396 458798
rect 580354 418296 580410 418305
rect 580354 418231 580410 418240
rect 580262 46336 580318 46345
rect 580262 46271 580318 46280
rect 580356 46232 580408 46238
rect 580356 46174 580408 46180
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 580368 19825 580396 46174
rect 580354 19816 580410 19825
rect 580354 19751 580410 19760
rect 575492 16546 575888 16574
rect 578252 16546 578648 16574
rect 574744 3868 574796 3874
rect 574744 3810 574796 3816
rect 572076 3392 572128 3398
rect 572076 3334 572128 3340
rect 572732 480 572760 3470
rect 574664 3454 575152 3482
rect 573916 3392 573968 3398
rect 573916 3334 573968 3340
rect 573928 480 573956 3334
rect 575124 480 575152 3454
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 567998 -960 568110 326
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 575860 354 575888 16546
rect 577412 3868 577464 3874
rect 577412 3810 577464 3816
rect 577424 480 577452 3810
rect 578620 480 578648 16546
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 581000 3596 581052 3602
rect 581000 3538 581052 3544
rect 581012 480 581040 3538
rect 582196 3460 582248 3466
rect 582196 3402 582248 3408
rect 582208 480 582236 3402
rect 583390 3360 583446 3369
rect 583390 3295 583446 3304
rect 583404 480 583432 3295
rect 576278 354 576390 480
rect 575860 326 576390 354
rect 576278 -960 576390 326
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3330 619112 3386 619168
rect 3330 606056 3386 606112
rect 3054 566888 3110 566944
rect 3330 553832 3386 553888
rect 3330 514820 3386 514856
rect 3330 514800 3332 514820
rect 3332 514800 3384 514820
rect 3384 514800 3386 514820
rect 3238 501744 3294 501800
rect 3514 671200 3570 671256
rect 3514 658144 3570 658200
rect 3514 632032 3570 632088
rect 3606 579944 3662 580000
rect 3698 527856 3754 527912
rect 3882 475632 3938 475688
rect 3514 462576 3570 462632
rect 3422 460128 3478 460184
rect 3514 449520 3570 449576
rect 3422 423544 3478 423600
rect 3422 410488 3478 410544
rect 3238 397432 3294 397488
rect 3238 371320 3294 371376
rect 3330 358400 3386 358456
rect 3146 345344 3202 345400
rect 3422 337320 3478 337376
rect 2778 306212 2780 306232
rect 2780 306212 2832 306232
rect 2832 306212 2834 306232
rect 2778 306176 2834 306212
rect 3054 293120 3110 293176
rect 3146 254088 3202 254144
rect 3330 214920 3386 214976
rect 3054 201864 3110 201920
rect 3238 162832 3294 162888
rect 4894 331744 4950 331800
rect 3514 319232 3570 319288
rect 3514 267144 3570 267200
rect 3514 241032 3570 241088
rect 3514 188808 3570 188864
rect 3422 136720 3478 136776
rect 3146 110608 3202 110664
rect 3422 84632 3478 84688
rect 3422 71576 3478 71632
rect 3422 32408 3478 32464
rect 3422 19352 3478 19408
rect 3514 6432 3570 6488
rect 5262 3304 5318 3360
rect 14554 330384 14610 330440
rect 90362 329024 90418 329080
rect 349158 460128 349214 460184
rect 244738 457408 244794 457464
rect 248970 457408 249026 457464
rect 252374 457408 252430 457464
rect 253662 457408 253718 457464
rect 258814 457408 258870 457464
rect 261942 457408 261998 457464
rect 263322 457408 263378 457464
rect 268198 457408 268254 457464
rect 271326 457408 271382 457464
rect 272890 457408 272946 457464
rect 385314 457408 385370 457464
rect 389638 457408 389694 457464
rect 394238 457408 394294 457464
rect 397550 457408 397606 457464
rect 398930 457408 398986 457464
rect 402058 457408 402114 457464
rect 403622 457408 403678 457464
rect 406750 457408 406806 457464
rect 408774 457408 408830 457464
rect 246302 338000 246358 338056
rect 250442 334056 250498 334112
rect 258170 3304 258226 3360
rect 282182 335960 282238 336016
rect 400862 338000 400918 338056
rect 392030 3304 392086 3360
rect 395434 334600 395490 334656
rect 396814 333240 396870 333296
rect 405002 327664 405058 327720
rect 407854 326304 407910 326360
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670656 580226 670712
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 432602 337456 432658 337512
rect 554042 164872 554098 164928
rect 580170 458088 580226 458144
rect 579618 431568 579674 431624
rect 579618 404912 579674 404968
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 580170 351872 580226 351928
rect 579894 325216 579950 325272
rect 580170 312024 580226 312080
rect 579618 298696 579674 298752
rect 579894 272176 579950 272232
rect 579802 258848 579858 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 580170 232328 580226 232384
rect 579894 219000 579950 219056
rect 580170 205672 580226 205728
rect 580170 192480 580226 192536
rect 579986 179152 580042 179208
rect 580170 165824 580226 165880
rect 579802 152632 579858 152688
rect 580170 125976 580226 126032
rect 580170 112784 580226 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 579986 72936 580042 72992
rect 580170 59608 580226 59664
rect 580354 418240 580410 418296
rect 580262 46280 580318 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 580354 19760 580410 19816
rect 580170 6568 580226 6624
rect 583390 3304 583446 3360
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3509 632090 3575 632093
rect -960 632088 3575 632090
rect -960 632032 3514 632088
rect 3570 632032 3575 632088
rect -960 632030 3575 632032
rect -960 631940 480 632030
rect 3509 632027 3575 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3325 619170 3391 619173
rect -960 619168 3391 619170
rect -960 619112 3330 619168
rect 3386 619112 3391 619168
rect -960 619110 3391 619112
rect -960 619020 480 619110
rect 3325 619107 3391 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3325 606114 3391 606117
rect -960 606112 3391 606114
rect -960 606056 3330 606112
rect 3386 606056 3391 606112
rect -960 606054 3391 606056
rect -960 605964 480 606054
rect 3325 606051 3391 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3601 580002 3667 580005
rect -960 580000 3667 580002
rect -960 579944 3606 580000
rect 3662 579944 3667 580000
rect -960 579942 3667 579944
rect -960 579852 480 579942
rect 3601 579939 3667 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3049 566946 3115 566949
rect -960 566944 3115 566946
rect -960 566888 3054 566944
rect 3110 566888 3115 566944
rect -960 566886 3115 566888
rect -960 566796 480 566886
rect 3049 566883 3115 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3693 527914 3759 527917
rect -960 527912 3759 527914
rect -960 527856 3698 527912
rect 3754 527856 3759 527912
rect -960 527854 3759 527856
rect -960 527764 480 527854
rect 3693 527851 3759 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3325 514858 3391 514861
rect -960 514856 3391 514858
rect -960 514800 3330 514856
rect 3386 514800 3391 514856
rect -960 514798 3391 514800
rect -960 514708 480 514798
rect 3325 514795 3391 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3233 501802 3299 501805
rect -960 501800 3299 501802
rect -960 501744 3238 501800
rect 3294 501744 3299 501800
rect -960 501742 3299 501744
rect -960 501652 480 501742
rect 3233 501739 3299 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3877 475690 3943 475693
rect -960 475688 3943 475690
rect -960 475632 3882 475688
rect 3938 475632 3943 475688
rect -960 475630 3943 475632
rect -960 475540 480 475630
rect 3877 475627 3943 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 3417 460186 3483 460189
rect 349153 460186 349219 460189
rect 3417 460184 349219 460186
rect 3417 460128 3422 460184
rect 3478 460128 349158 460184
rect 349214 460128 349219 460184
rect 3417 460126 349219 460128
rect 3417 460123 3483 460126
rect 349153 460123 349219 460126
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 244733 457466 244799 457469
rect 248965 457468 249031 457469
rect 252369 457468 252435 457469
rect 253657 457468 253723 457469
rect 245510 457466 245516 457468
rect 244733 457464 245516 457466
rect 244733 457408 244738 457464
rect 244794 457408 245516 457464
rect 244733 457406 245516 457408
rect 244733 457403 244799 457406
rect 245510 457404 245516 457406
rect 245580 457404 245586 457468
rect 248965 457464 249012 457468
rect 249076 457466 249082 457468
rect 252318 457466 252324 457468
rect 248965 457408 248970 457464
rect 248965 457404 249012 457408
rect 249076 457406 249122 457466
rect 252278 457406 252324 457466
rect 252388 457464 252435 457468
rect 253606 457466 253612 457468
rect 252430 457408 252435 457464
rect 249076 457404 249082 457406
rect 252318 457404 252324 457406
rect 252388 457404 252435 457408
rect 253566 457406 253612 457466
rect 253676 457464 253723 457468
rect 253718 457408 253723 457464
rect 253606 457404 253612 457406
rect 253676 457404 253723 457408
rect 248965 457403 249031 457404
rect 252369 457403 252435 457404
rect 253657 457403 253723 457404
rect 258809 457466 258875 457469
rect 259310 457466 259316 457468
rect 258809 457464 259316 457466
rect 258809 457408 258814 457464
rect 258870 457408 259316 457464
rect 258809 457406 259316 457408
rect 258809 457403 258875 457406
rect 259310 457404 259316 457406
rect 259380 457404 259386 457468
rect 261937 457466 262003 457469
rect 263317 457468 263383 457469
rect 262070 457466 262076 457468
rect 261937 457464 262076 457466
rect 261937 457408 261942 457464
rect 261998 457408 262076 457464
rect 261937 457406 262076 457408
rect 261937 457403 262003 457406
rect 262070 457404 262076 457406
rect 262140 457404 262146 457468
rect 263317 457464 263364 457468
rect 263428 457466 263434 457468
rect 268193 457466 268259 457469
rect 268878 457466 268884 457468
rect 263317 457408 263322 457464
rect 263317 457404 263364 457408
rect 263428 457406 263474 457466
rect 268193 457464 268884 457466
rect 268193 457408 268198 457464
rect 268254 457408 268884 457464
rect 268193 457406 268884 457408
rect 263428 457404 263434 457406
rect 263317 457403 263383 457404
rect 268193 457403 268259 457406
rect 268878 457404 268884 457406
rect 268948 457404 268954 457468
rect 271321 457466 271387 457469
rect 271638 457466 271644 457468
rect 271321 457464 271644 457466
rect 271321 457408 271326 457464
rect 271382 457408 271644 457464
rect 271321 457406 271644 457408
rect 271321 457403 271387 457406
rect 271638 457404 271644 457406
rect 271708 457404 271714 457468
rect 272885 457466 272951 457469
rect 273110 457466 273116 457468
rect 272885 457464 273116 457466
rect 272885 457408 272890 457464
rect 272946 457408 273116 457464
rect 272885 457406 273116 457408
rect 272885 457403 272951 457406
rect 273110 457404 273116 457406
rect 273180 457404 273186 457468
rect 385166 457404 385172 457468
rect 385236 457466 385242 457468
rect 385309 457466 385375 457469
rect 389633 457468 389699 457469
rect 389582 457466 389588 457468
rect 385236 457464 385375 457466
rect 385236 457408 385314 457464
rect 385370 457408 385375 457464
rect 385236 457406 385375 457408
rect 389542 457406 389588 457466
rect 389652 457464 389699 457468
rect 389694 457408 389699 457464
rect 385236 457404 385242 457406
rect 385309 457403 385375 457406
rect 389582 457404 389588 457406
rect 389652 457404 389699 457408
rect 393998 457404 394004 457468
rect 394068 457466 394074 457468
rect 394233 457466 394299 457469
rect 397545 457468 397611 457469
rect 397494 457466 397500 457468
rect 394068 457464 394299 457466
rect 394068 457408 394238 457464
rect 394294 457408 394299 457464
rect 394068 457406 394299 457408
rect 397454 457406 397500 457466
rect 397564 457464 397611 457468
rect 397606 457408 397611 457464
rect 394068 457404 394074 457406
rect 389633 457403 389699 457404
rect 394233 457403 394299 457406
rect 397494 457404 397500 457406
rect 397564 457404 397611 457408
rect 398782 457404 398788 457468
rect 398852 457466 398858 457468
rect 398925 457466 398991 457469
rect 398852 457464 398991 457466
rect 398852 457408 398930 457464
rect 398986 457408 398991 457464
rect 398852 457406 398991 457408
rect 398852 457404 398858 457406
rect 397545 457403 397611 457404
rect 398925 457403 398991 457406
rect 401542 457404 401548 457468
rect 401612 457466 401618 457468
rect 402053 457466 402119 457469
rect 401612 457464 402119 457466
rect 401612 457408 402058 457464
rect 402114 457408 402119 457464
rect 401612 457406 402119 457408
rect 401612 457404 401618 457406
rect 402053 457403 402119 457406
rect 403014 457404 403020 457468
rect 403084 457466 403090 457468
rect 403617 457466 403683 457469
rect 403084 457464 403683 457466
rect 403084 457408 403622 457464
rect 403678 457408 403683 457464
rect 403084 457406 403683 457408
rect 403084 457404 403090 457406
rect 403617 457403 403683 457406
rect 405774 457404 405780 457468
rect 405844 457466 405850 457468
rect 406745 457466 406811 457469
rect 408769 457468 408835 457469
rect 408718 457466 408724 457468
rect 405844 457464 406811 457466
rect 405844 457408 406750 457464
rect 406806 457408 406811 457464
rect 405844 457406 406811 457408
rect 408678 457406 408724 457466
rect 408788 457464 408835 457468
rect 408830 457408 408835 457464
rect 405844 457404 405850 457406
rect 406745 457403 406811 457406
rect 408718 457404 408724 457406
rect 408788 457404 408835 457408
rect 408769 457403 408835 457404
rect -960 449578 480 449668
rect 3509 449578 3575 449581
rect -960 449576 3575 449578
rect -960 449520 3514 449576
rect 3570 449520 3575 449576
rect -960 449518 3575 449520
rect -960 449428 480 449518
rect 3509 449515 3575 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 579613 431626 579679 431629
rect 583520 431626 584960 431716
rect 579613 431624 584960 431626
rect 579613 431568 579618 431624
rect 579674 431568 584960 431624
rect 579613 431566 584960 431568
rect 579613 431563 579679 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 580349 418298 580415 418301
rect 583520 418298 584960 418388
rect 580349 418296 584960 418298
rect 580349 418240 580354 418296
rect 580410 418240 584960 418296
rect 580349 418238 584960 418240
rect 580349 418235 580415 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3417 410546 3483 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect -960 410486 3483 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 579613 404970 579679 404973
rect 583520 404970 584960 405060
rect 579613 404968 584960 404970
rect 579613 404912 579618 404968
rect 579674 404912 584960 404968
rect 579613 404910 584960 404912
rect 579613 404907 579679 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3233 397490 3299 397493
rect -960 397488 3299 397490
rect -960 397432 3238 397488
rect 3294 397432 3299 397488
rect -960 397430 3299 397432
rect -960 397340 480 397430
rect 3233 397427 3299 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3233 371378 3299 371381
rect -960 371376 3299 371378
rect -960 371320 3238 371376
rect 3294 371320 3299 371376
rect -960 371318 3299 371320
rect -960 371228 480 371318
rect 3233 371315 3299 371318
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3141 345402 3207 345405
rect -960 345400 3207 345402
rect -960 345344 3146 345400
rect 3202 345344 3207 345400
rect -960 345342 3207 345344
rect -960 345252 480 345342
rect 3141 345339 3207 345342
rect 583520 338452 584960 338692
rect 245510 337996 245516 338060
rect 245580 338058 245586 338060
rect 246297 338058 246363 338061
rect 245580 338056 246363 338058
rect 245580 338000 246302 338056
rect 246358 338000 246363 338056
rect 245580 337998 246363 338000
rect 245580 337996 245586 337998
rect 246297 337995 246363 337998
rect 400857 338058 400923 338061
rect 401542 338058 401548 338060
rect 400857 338056 401548 338058
rect 400857 338000 400862 338056
rect 400918 338000 401548 338056
rect 400857 337998 401548 338000
rect 400857 337995 400923 337998
rect 401542 337996 401548 337998
rect 401612 337996 401618 338060
rect 263358 337452 263364 337516
rect 263428 337514 263434 337516
rect 432597 337514 432663 337517
rect 263428 337512 432663 337514
rect 263428 337456 432602 337512
rect 432658 337456 432663 337512
rect 263428 337454 432663 337456
rect 263428 337452 263434 337454
rect 432597 337451 432663 337454
rect 3417 337378 3483 337381
rect 397494 337378 397500 337380
rect 3417 337376 397500 337378
rect 3417 337320 3422 337376
rect 3478 337320 397500 337376
rect 3417 337318 397500 337320
rect 3417 337315 3483 337318
rect 397494 337316 397500 337318
rect 397564 337316 397570 337380
rect 273110 335956 273116 336020
rect 273180 336018 273186 336020
rect 282177 336018 282243 336021
rect 273180 336016 282243 336018
rect 273180 335960 282182 336016
rect 282238 335960 282243 336016
rect 273180 335958 282243 335960
rect 273180 335956 273186 335958
rect 282177 335955 282243 335958
rect 262070 334596 262076 334660
rect 262140 334658 262146 334660
rect 395429 334658 395495 334661
rect 262140 334656 395495 334658
rect 262140 334600 395434 334656
rect 395490 334600 395495 334656
rect 262140 334598 395495 334600
rect 262140 334596 262146 334598
rect 395429 334595 395495 334598
rect 249006 334052 249012 334116
rect 249076 334114 249082 334116
rect 250437 334114 250503 334117
rect 249076 334112 250503 334114
rect 249076 334056 250442 334112
rect 250498 334056 250503 334112
rect 249076 334054 250503 334056
rect 249076 334052 249082 334054
rect 250437 334051 250503 334054
rect 271638 333236 271644 333300
rect 271708 333298 271714 333300
rect 396809 333298 396875 333301
rect 271708 333296 396875 333298
rect 271708 333240 396814 333296
rect 396870 333240 396875 333296
rect 271708 333238 396875 333240
rect 271708 333236 271714 333238
rect 396809 333235 396875 333238
rect -960 332196 480 332436
rect 4889 331802 4955 331805
rect 385166 331802 385172 331804
rect 4889 331800 385172 331802
rect 4889 331744 4894 331800
rect 4950 331744 385172 331800
rect 4889 331742 385172 331744
rect 4889 331739 4955 331742
rect 385166 331740 385172 331742
rect 385236 331740 385242 331804
rect 14549 330442 14615 330445
rect 389582 330442 389588 330444
rect 14549 330440 389588 330442
rect 14549 330384 14554 330440
rect 14610 330384 389588 330440
rect 14549 330382 389588 330384
rect 14549 330379 14615 330382
rect 389582 330380 389588 330382
rect 389652 330380 389658 330444
rect 90357 329082 90423 329085
rect 393998 329082 394004 329084
rect 90357 329080 394004 329082
rect 90357 329024 90362 329080
rect 90418 329024 394004 329080
rect 90357 329022 394004 329024
rect 90357 329019 90423 329022
rect 393998 329020 394004 329022
rect 394068 329020 394074 329084
rect 259310 327660 259316 327724
rect 259380 327722 259386 327724
rect 404997 327722 405063 327725
rect 259380 327720 405063 327722
rect 259380 327664 405002 327720
rect 405058 327664 405063 327720
rect 259380 327662 405063 327664
rect 259380 327660 259386 327662
rect 404997 327659 405063 327662
rect 268878 326300 268884 326364
rect 268948 326362 268954 326364
rect 407849 326362 407915 326365
rect 268948 326360 407915 326362
rect 268948 326304 407854 326360
rect 407910 326304 407915 326360
rect 268948 326302 407915 326304
rect 268948 326300 268954 326302
rect 407849 326299 407915 326302
rect 579889 325274 579955 325277
rect 583520 325274 584960 325364
rect 579889 325272 584960 325274
rect 579889 325216 579894 325272
rect 579950 325216 584960 325272
rect 579889 325214 584960 325216
rect 579889 325211 579955 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3509 319290 3575 319293
rect -960 319288 3575 319290
rect -960 319232 3514 319288
rect 3570 319232 3575 319288
rect -960 319230 3575 319232
rect -960 319140 480 319230
rect 3509 319227 3575 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 2773 306234 2839 306237
rect -960 306232 2839 306234
rect -960 306176 2778 306232
rect 2834 306176 2839 306232
rect -960 306174 2839 306176
rect -960 306084 480 306174
rect 2773 306171 2839 306174
rect 579613 298754 579679 298757
rect 583520 298754 584960 298844
rect 579613 298752 584960 298754
rect 579613 298696 579618 298752
rect 579674 298696 584960 298752
rect 579613 298694 584960 298696
rect 579613 298691 579679 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3049 293178 3115 293181
rect -960 293176 3115 293178
rect -960 293120 3054 293176
rect 3110 293120 3115 293176
rect -960 293118 3115 293120
rect -960 293028 480 293118
rect 3049 293115 3115 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 579889 272234 579955 272237
rect 583520 272234 584960 272324
rect 579889 272232 584960 272234
rect 579889 272176 579894 272232
rect 579950 272176 584960 272232
rect 579889 272174 584960 272176
rect 579889 272171 579955 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3509 267202 3575 267205
rect -960 267200 3575 267202
rect -960 267144 3514 267200
rect 3570 267144 3575 267200
rect -960 267142 3575 267144
rect -960 267052 480 267142
rect 3509 267139 3575 267142
rect 579797 258906 579863 258909
rect 583520 258906 584960 258996
rect 579797 258904 584960 258906
rect 579797 258848 579802 258904
rect 579858 258848 584960 258904
rect 579797 258846 584960 258848
rect 579797 258843 579863 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 579889 219058 579955 219061
rect 583520 219058 584960 219148
rect 579889 219056 584960 219058
rect 579889 219000 579894 219056
rect 579950 219000 584960 219056
rect 579889 218998 584960 219000
rect 579889 218995 579955 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3049 201922 3115 201925
rect -960 201920 3115 201922
rect -960 201864 3054 201920
rect 3110 201864 3115 201920
rect -960 201862 3115 201864
rect -960 201772 480 201862
rect 3049 201859 3115 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 579981 179210 580047 179213
rect 583520 179210 584960 179300
rect 579981 179208 584960 179210
rect 579981 179152 579986 179208
rect 580042 179152 584960 179208
rect 579981 179150 584960 179152
rect 579981 179147 580047 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect 252318 164868 252324 164932
rect 252388 164930 252394 164932
rect 554037 164930 554103 164933
rect 252388 164928 554103 164930
rect 252388 164872 554042 164928
rect 554098 164872 554103 164928
rect 252388 164870 554103 164872
rect 252388 164868 252394 164870
rect 554037 164867 554103 164870
rect -960 162890 480 162980
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 579797 152690 579863 152693
rect 583520 152690 584960 152780
rect 579797 152688 584960 152690
rect 579797 152632 579802 152688
rect 579858 152632 584960 152688
rect 579797 152630 584960 152632
rect 579797 152627 579863 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect -960 149774 674 149834
rect -960 149698 480 149774
rect 614 149698 674 149774
rect -960 149684 674 149698
rect 246 149638 674 149684
rect 246 149154 306 149638
rect 398782 149154 398788 149156
rect 246 149094 398788 149154
rect 398782 149092 398788 149094
rect 398852 149092 398858 149156
rect 583520 139362 584960 139452
rect 583342 139302 584960 139362
rect 583342 139226 583402 139302
rect 583520 139226 584960 139302
rect 583342 139212 584960 139226
rect 583342 139166 583586 139212
rect 253606 138076 253612 138140
rect 253676 138138 253682 138140
rect 583526 138138 583586 139166
rect 253676 138078 583586 138138
rect 253676 138076 253682 138078
rect -960 136778 480 136868
rect 3417 136778 3483 136781
rect -960 136776 3483 136778
rect -960 136720 3422 136776
rect 3478 136720 3483 136776
rect -960 136718 3483 136720
rect -960 136628 480 136718
rect 3417 136715 3483 136718
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 580165 112842 580231 112845
rect 583520 112842 584960 112932
rect 580165 112840 584960 112842
rect 580165 112784 580170 112840
rect 580226 112784 584960 112840
rect 580165 112782 584960 112784
rect 580165 112779 580231 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect -960 97550 674 97610
rect -960 97474 480 97550
rect 614 97474 674 97550
rect -960 97460 674 97474
rect 246 97414 674 97460
rect 246 96930 306 97414
rect 246 96870 6930 96930
rect 6870 96658 6930 96870
rect 403014 96658 403020 96660
rect 6870 96598 403020 96658
rect 403014 96596 403020 96598
rect 403084 96596 403090 96660
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3417 84690 3483 84693
rect -960 84688 3483 84690
rect -960 84632 3422 84688
rect 3478 84632 3483 84688
rect -960 84630 3483 84632
rect -960 84540 480 84630
rect 3417 84627 3483 84630
rect 579981 72994 580047 72997
rect 583520 72994 584960 73084
rect 579981 72992 584960 72994
rect 579981 72936 579986 72992
rect 580042 72936 584960 72992
rect 579981 72934 584960 72936
rect 579981 72931 580047 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect -960 58518 674 58578
rect -960 58442 480 58518
rect 614 58442 674 58518
rect -960 58428 674 58442
rect 246 58382 674 58428
rect 246 58034 306 58382
rect 408718 58034 408724 58036
rect 246 57974 408724 58034
rect 408718 57972 408724 57974
rect 408788 57972 408794 58036
rect 580257 46338 580323 46341
rect 583520 46338 584960 46428
rect 580257 46336 584960 46338
rect 580257 46280 580262 46336
rect 580318 46280 584960 46336
rect 580257 46278 584960 46280
rect 580257 46275 580323 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect -960 45462 674 45522
rect -960 45386 480 45462
rect 614 45386 674 45462
rect -960 45372 674 45386
rect 246 45326 674 45372
rect 246 44842 306 45326
rect 246 44782 6930 44842
rect 6870 44298 6930 44782
rect 405774 44298 405780 44300
rect 6870 44238 405780 44298
rect 405774 44236 405780 44238
rect 405844 44236 405850 44300
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3417 32466 3483 32469
rect -960 32464 3483 32466
rect -960 32408 3422 32464
rect 3478 32408 3483 32464
rect -960 32406 3483 32408
rect -960 32316 480 32406
rect 3417 32403 3483 32406
rect 580349 19818 580415 19821
rect 583520 19818 584960 19908
rect 580349 19816 584960 19818
rect 580349 19760 580354 19816
rect 580410 19760 584960 19816
rect 580349 19758 584960 19760
rect 580349 19755 580415 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3509 6490 3575 6493
rect -960 6488 3575 6490
rect -960 6432 3514 6488
rect 3570 6432 3575 6488
rect 583520 6476 584960 6566
rect -960 6430 3575 6432
rect -960 6340 480 6430
rect 3509 6427 3575 6430
rect 5257 3362 5323 3365
rect 258165 3362 258231 3365
rect 5257 3360 258231 3362
rect 5257 3304 5262 3360
rect 5318 3304 258170 3360
rect 258226 3304 258231 3360
rect 5257 3302 258231 3304
rect 5257 3299 5323 3302
rect 258165 3299 258231 3302
rect 392025 3362 392091 3365
rect 583385 3362 583451 3365
rect 392025 3360 583451 3362
rect 392025 3304 392030 3360
rect 392086 3304 583390 3360
rect 583446 3304 583451 3360
rect 392025 3302 583451 3304
rect 392025 3299 392091 3302
rect 583385 3299 583451 3302
<< via3 >>
rect 245516 457404 245580 457468
rect 249012 457464 249076 457468
rect 249012 457408 249026 457464
rect 249026 457408 249076 457464
rect 249012 457404 249076 457408
rect 252324 457464 252388 457468
rect 252324 457408 252374 457464
rect 252374 457408 252388 457464
rect 252324 457404 252388 457408
rect 253612 457464 253676 457468
rect 253612 457408 253662 457464
rect 253662 457408 253676 457464
rect 253612 457404 253676 457408
rect 259316 457404 259380 457468
rect 262076 457404 262140 457468
rect 263364 457464 263428 457468
rect 263364 457408 263378 457464
rect 263378 457408 263428 457464
rect 263364 457404 263428 457408
rect 268884 457404 268948 457468
rect 271644 457404 271708 457468
rect 273116 457404 273180 457468
rect 385172 457404 385236 457468
rect 389588 457464 389652 457468
rect 389588 457408 389638 457464
rect 389638 457408 389652 457464
rect 389588 457404 389652 457408
rect 394004 457404 394068 457468
rect 397500 457464 397564 457468
rect 397500 457408 397550 457464
rect 397550 457408 397564 457464
rect 397500 457404 397564 457408
rect 398788 457404 398852 457468
rect 401548 457404 401612 457468
rect 403020 457404 403084 457468
rect 405780 457404 405844 457468
rect 408724 457464 408788 457468
rect 408724 457408 408774 457464
rect 408774 457408 408788 457464
rect 408724 457404 408788 457408
rect 245516 337996 245580 338060
rect 401548 337996 401612 338060
rect 263364 337452 263428 337516
rect 397500 337316 397564 337380
rect 273116 335956 273180 336020
rect 262076 334596 262140 334660
rect 249012 334052 249076 334116
rect 271644 333236 271708 333300
rect 385172 331740 385236 331804
rect 389588 330380 389652 330444
rect 394004 329020 394068 329084
rect 259316 327660 259380 327724
rect 268884 326300 268948 326364
rect 252324 164868 252388 164932
rect 398788 149092 398852 149156
rect 253612 138076 253676 138140
rect 403020 96596 403084 96660
rect 408724 57972 408788 58036
rect 405780 44236 405844 44300
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 205954 96914 241398
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 210454 101414 245898
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100794 174454 101414 209898
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 214954 105914 250398
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 223954 114914 259398
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114294 115954 114914 151398
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 228454 119414 263898
rect 118794 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 119414 228454
rect 118794 228134 119414 228218
rect 118794 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 119414 228134
rect 118794 192454 119414 227898
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 120454 119414 155898
rect 118794 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 119414 120454
rect 118794 120134 119414 120218
rect 118794 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 119414 120134
rect 118794 84454 119414 119898
rect 118794 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 119414 84454
rect 118794 84134 119414 84218
rect 118794 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 119414 84134
rect 118794 48454 119414 83898
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 232954 123914 268398
rect 123294 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 123914 232954
rect 123294 232634 123914 232718
rect 123294 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 123914 232634
rect 123294 196954 123914 232398
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 124954 123914 160398
rect 123294 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 123914 124954
rect 123294 124634 123914 124718
rect 123294 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 123914 124634
rect 123294 88954 123914 124398
rect 123294 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 123914 88954
rect 123294 88634 123914 88718
rect 123294 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 123914 88634
rect 123294 52954 123914 88398
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 241954 132914 277398
rect 132294 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 132914 241954
rect 132294 241634 132914 241718
rect 132294 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 132914 241634
rect 132294 205954 132914 241398
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 132294 169954 132914 205398
rect 132294 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 132914 169954
rect 132294 169634 132914 169718
rect 132294 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 132914 169634
rect 132294 133954 132914 169398
rect 132294 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 132914 133954
rect 132294 133634 132914 133718
rect 132294 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 132914 133634
rect 132294 97954 132914 133398
rect 132294 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 132914 97954
rect 132294 97634 132914 97718
rect 132294 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 132914 97634
rect 132294 61954 132914 97398
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 246454 137414 281898
rect 136794 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 137414 246454
rect 136794 246134 137414 246218
rect 136794 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 137414 246134
rect 136794 210454 137414 245898
rect 136794 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 137414 210454
rect 136794 210134 137414 210218
rect 136794 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 137414 210134
rect 136794 174454 137414 209898
rect 136794 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 137414 174454
rect 136794 174134 137414 174218
rect 136794 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 137414 174134
rect 136794 138454 137414 173898
rect 136794 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 137414 138454
rect 136794 138134 137414 138218
rect 136794 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 137414 138134
rect 136794 102454 137414 137898
rect 136794 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 137414 102454
rect 136794 102134 137414 102218
rect 136794 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 137414 102134
rect 136794 66454 137414 101898
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 214954 141914 250398
rect 141294 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 141914 214954
rect 141294 214634 141914 214718
rect 141294 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 141914 214634
rect 141294 178954 141914 214398
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 141294 142954 141914 178398
rect 141294 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 141914 142954
rect 141294 142634 141914 142718
rect 141294 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 141914 142634
rect 141294 106954 141914 142398
rect 141294 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 141914 106954
rect 141294 106634 141914 106718
rect 141294 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 141914 106634
rect 141294 70954 141914 106398
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 223954 150914 259398
rect 150294 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 150914 223954
rect 150294 223634 150914 223718
rect 150294 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 150914 223634
rect 150294 187954 150914 223398
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 150294 151954 150914 187398
rect 150294 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 150914 151954
rect 150294 151634 150914 151718
rect 150294 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 150914 151634
rect 150294 115954 150914 151398
rect 150294 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 150914 115954
rect 150294 115634 150914 115718
rect 150294 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 150914 115634
rect 150294 79954 150914 115398
rect 150294 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 150914 79954
rect 150294 79634 150914 79718
rect 150294 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 150914 79634
rect 150294 43954 150914 79398
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 228454 155414 263898
rect 154794 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 155414 228454
rect 154794 228134 155414 228218
rect 154794 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 155414 228134
rect 154794 192454 155414 227898
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154794 156454 155414 191898
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154794 120454 155414 155898
rect 154794 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 155414 120454
rect 154794 120134 155414 120218
rect 154794 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 155414 120134
rect 154794 84454 155414 119898
rect 154794 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 155414 84454
rect 154794 84134 155414 84218
rect 154794 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 155414 84134
rect 154794 48454 155414 83898
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 232954 159914 268398
rect 159294 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 159914 232954
rect 159294 232634 159914 232718
rect 159294 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 159914 232634
rect 159294 196954 159914 232398
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 159294 160954 159914 196398
rect 159294 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 159914 160954
rect 159294 160634 159914 160718
rect 159294 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 159914 160634
rect 159294 124954 159914 160398
rect 159294 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 159914 124954
rect 159294 124634 159914 124718
rect 159294 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 159914 124634
rect 159294 88954 159914 124398
rect 159294 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 159914 88954
rect 159294 88634 159914 88718
rect 159294 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 159914 88634
rect 159294 52954 159914 88398
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 241954 168914 277398
rect 168294 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 168914 241954
rect 168294 241634 168914 241718
rect 168294 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 168914 241634
rect 168294 205954 168914 241398
rect 168294 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 168914 205954
rect 168294 205634 168914 205718
rect 168294 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 168914 205634
rect 168294 169954 168914 205398
rect 168294 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 168914 169954
rect 168294 169634 168914 169718
rect 168294 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 168914 169634
rect 168294 133954 168914 169398
rect 168294 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 168914 133954
rect 168294 133634 168914 133718
rect 168294 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 168914 133634
rect 168294 97954 168914 133398
rect 168294 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 168914 97954
rect 168294 97634 168914 97718
rect 168294 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 168914 97634
rect 168294 61954 168914 97398
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 246454 173414 281898
rect 172794 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 173414 246454
rect 172794 246134 173414 246218
rect 172794 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 173414 246134
rect 172794 210454 173414 245898
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 172794 138454 173414 173898
rect 172794 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 173414 138454
rect 172794 138134 173414 138218
rect 172794 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 173414 138134
rect 172794 102454 173414 137898
rect 172794 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 173414 102454
rect 172794 102134 173414 102218
rect 172794 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 173414 102134
rect 172794 66454 173414 101898
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 214954 177914 250398
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 106954 177914 142398
rect 177294 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 177914 106954
rect 177294 106634 177914 106718
rect 177294 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 177914 106634
rect 177294 70954 177914 106398
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 223954 186914 259398
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 186294 79954 186914 115398
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 228454 191414 263898
rect 190794 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 191414 228454
rect 190794 228134 191414 228218
rect 190794 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 191414 228134
rect 190794 192454 191414 227898
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 232954 195914 268398
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 205954 204914 241398
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 210454 209414 245898
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 214954 213914 250398
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 223954 222914 259398
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 228454 227414 263898
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 226794 192454 227414 227898
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 460000 236414 488898
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 460000 240914 493398
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 460000 245414 461898
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 460000 249914 466398
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 460000 254414 470898
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 460000 258914 475398
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 460000 263414 479898
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 460000 267914 484398
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 460000 272414 488898
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 460000 276914 493398
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 460000 281414 461898
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 460000 285914 466398
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 460000 290414 470898
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 460000 294914 475398
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 460000 299414 479898
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 460000 303914 484398
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 460000 308414 488898
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 460000 312914 493398
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 460000 317414 461898
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 460000 321914 466398
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 460000 326414 470898
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 460000 330914 475398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 460000 335414 479898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 460000 339914 484398
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 460000 344414 488898
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 460000 348914 493398
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 460000 353414 461898
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 460000 357914 466398
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 460000 362414 470898
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 460000 366914 475398
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 460000 371414 479898
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 460000 375914 484398
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 460000 380414 488898
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 460000 384914 493398
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 460000 389414 461898
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 460000 393914 466398
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 460000 398414 470898
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 460000 402914 475398
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 460000 407414 479898
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 460000 411914 484398
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 460000 416414 488898
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 245515 457468 245581 457469
rect 245515 457404 245516 457468
rect 245580 457404 245581 457468
rect 245515 457403 245581 457404
rect 249011 457468 249077 457469
rect 249011 457404 249012 457468
rect 249076 457404 249077 457468
rect 249011 457403 249077 457404
rect 252323 457468 252389 457469
rect 252323 457404 252324 457468
rect 252388 457404 252389 457468
rect 252323 457403 252389 457404
rect 253611 457468 253677 457469
rect 253611 457404 253612 457468
rect 253676 457404 253677 457468
rect 253611 457403 253677 457404
rect 259315 457468 259381 457469
rect 259315 457404 259316 457468
rect 259380 457404 259381 457468
rect 259315 457403 259381 457404
rect 262075 457468 262141 457469
rect 262075 457404 262076 457468
rect 262140 457404 262141 457468
rect 262075 457403 262141 457404
rect 263363 457468 263429 457469
rect 263363 457404 263364 457468
rect 263428 457404 263429 457468
rect 263363 457403 263429 457404
rect 268883 457468 268949 457469
rect 268883 457404 268884 457468
rect 268948 457404 268949 457468
rect 268883 457403 268949 457404
rect 271643 457468 271709 457469
rect 271643 457404 271644 457468
rect 271708 457404 271709 457468
rect 271643 457403 271709 457404
rect 273115 457468 273181 457469
rect 273115 457404 273116 457468
rect 273180 457404 273181 457468
rect 273115 457403 273181 457404
rect 385171 457468 385237 457469
rect 385171 457404 385172 457468
rect 385236 457404 385237 457468
rect 385171 457403 385237 457404
rect 389587 457468 389653 457469
rect 389587 457404 389588 457468
rect 389652 457404 389653 457468
rect 389587 457403 389653 457404
rect 394003 457468 394069 457469
rect 394003 457404 394004 457468
rect 394068 457404 394069 457468
rect 394003 457403 394069 457404
rect 397499 457468 397565 457469
rect 397499 457404 397500 457468
rect 397564 457404 397565 457468
rect 397499 457403 397565 457404
rect 398787 457468 398853 457469
rect 398787 457404 398788 457468
rect 398852 457404 398853 457468
rect 398787 457403 398853 457404
rect 401547 457468 401613 457469
rect 401547 457404 401548 457468
rect 401612 457404 401613 457468
rect 401547 457403 401613 457404
rect 403019 457468 403085 457469
rect 403019 457404 403020 457468
rect 403084 457404 403085 457468
rect 403019 457403 403085 457404
rect 405779 457468 405845 457469
rect 405779 457404 405780 457468
rect 405844 457404 405845 457468
rect 405779 457403 405845 457404
rect 408723 457468 408789 457469
rect 408723 457404 408724 457468
rect 408788 457404 408789 457468
rect 408723 457403 408789 457404
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 239208 435454 239528 435486
rect 239208 435218 239250 435454
rect 239486 435218 239528 435454
rect 239208 435134 239528 435218
rect 239208 434898 239250 435134
rect 239486 434898 239528 435134
rect 239208 434866 239528 434898
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 239208 399454 239528 399486
rect 239208 399218 239250 399454
rect 239486 399218 239528 399454
rect 239208 399134 239528 399218
rect 239208 398898 239250 399134
rect 239486 398898 239528 399134
rect 239208 398866 239528 398898
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 239208 363454 239528 363486
rect 239208 363218 239250 363454
rect 239486 363218 239528 363454
rect 239208 363134 239528 363218
rect 239208 362898 239250 363134
rect 239486 362898 239528 363134
rect 239208 362866 239528 362898
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 245518 338061 245578 457403
rect 245515 338060 245581 338061
rect 245515 337996 245516 338060
rect 245580 337996 245581 338060
rect 245515 337995 245581 337996
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 232954 231914 268398
rect 231294 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 231914 232954
rect 231294 232634 231914 232718
rect 231294 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 231914 232634
rect 231294 196954 231914 232398
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 309454 236414 336000
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 313954 240914 336000
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 241954 240914 277398
rect 240294 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 240914 241954
rect 240294 241634 240914 241718
rect 240294 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 240914 241634
rect 240294 205954 240914 241398
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 318454 245414 336000
rect 249014 334117 249074 457403
rect 249011 334116 249077 334117
rect 249011 334052 249012 334116
rect 249076 334052 249077 334116
rect 249011 334051 249077 334052
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 210454 245414 245898
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 322954 249914 336000
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 214954 249914 250398
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 252326 164933 252386 457403
rect 252323 164932 252389 164933
rect 252323 164868 252324 164932
rect 252388 164868 252389 164932
rect 252323 164867 252389 164868
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 253614 138141 253674 457403
rect 254568 439954 254888 439986
rect 254568 439718 254610 439954
rect 254846 439718 254888 439954
rect 254568 439634 254888 439718
rect 254568 439398 254610 439634
rect 254846 439398 254888 439634
rect 254568 439366 254888 439398
rect 254568 403954 254888 403986
rect 254568 403718 254610 403954
rect 254846 403718 254888 403954
rect 254568 403634 254888 403718
rect 254568 403398 254610 403634
rect 254846 403398 254888 403634
rect 254568 403366 254888 403398
rect 254568 367954 254888 367986
rect 254568 367718 254610 367954
rect 254846 367718 254888 367954
rect 254568 367634 254888 367718
rect 254568 367398 254610 367634
rect 254846 367398 254888 367634
rect 254568 367366 254888 367398
rect 253794 327454 254414 336000
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253611 138140 253677 138141
rect 253611 138076 253612 138140
rect 253676 138076 253677 138140
rect 253611 138075 253677 138076
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 331954 258914 336000
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 259318 327725 259378 457403
rect 262078 334661 262138 457403
rect 263366 337517 263426 457403
rect 263363 337516 263429 337517
rect 263363 337452 263364 337516
rect 263428 337452 263429 337516
rect 263363 337451 263429 337452
rect 262075 334660 262141 334661
rect 262075 334596 262076 334660
rect 262140 334596 262141 334660
rect 262075 334595 262141 334596
rect 259315 327724 259381 327725
rect 259315 327660 259316 327724
rect 259380 327660 259381 327724
rect 259315 327659 259381 327660
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 223954 258914 259398
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 300454 263414 336000
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 228454 263414 263898
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 262794 192454 263414 227898
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 304954 267914 336000
rect 268886 326365 268946 457403
rect 269928 435454 270248 435486
rect 269928 435218 269970 435454
rect 270206 435218 270248 435454
rect 269928 435134 270248 435218
rect 269928 434898 269970 435134
rect 270206 434898 270248 435134
rect 269928 434866 270248 434898
rect 269928 399454 270248 399486
rect 269928 399218 269970 399454
rect 270206 399218 270248 399454
rect 269928 399134 270248 399218
rect 269928 398898 269970 399134
rect 270206 398898 270248 399134
rect 269928 398866 270248 398898
rect 269928 363454 270248 363486
rect 269928 363218 269970 363454
rect 270206 363218 270248 363454
rect 269928 363134 270248 363218
rect 269928 362898 269970 363134
rect 270206 362898 270248 363134
rect 269928 362866 270248 362898
rect 271646 333301 271706 457403
rect 273118 336021 273178 457403
rect 285288 439954 285608 439986
rect 285288 439718 285330 439954
rect 285566 439718 285608 439954
rect 285288 439634 285608 439718
rect 285288 439398 285330 439634
rect 285566 439398 285608 439634
rect 285288 439366 285608 439398
rect 316008 439954 316328 439986
rect 316008 439718 316050 439954
rect 316286 439718 316328 439954
rect 316008 439634 316328 439718
rect 316008 439398 316050 439634
rect 316286 439398 316328 439634
rect 316008 439366 316328 439398
rect 346728 439954 347048 439986
rect 346728 439718 346770 439954
rect 347006 439718 347048 439954
rect 346728 439634 347048 439718
rect 346728 439398 346770 439634
rect 347006 439398 347048 439634
rect 346728 439366 347048 439398
rect 377448 439954 377768 439986
rect 377448 439718 377490 439954
rect 377726 439718 377768 439954
rect 377448 439634 377768 439718
rect 377448 439398 377490 439634
rect 377726 439398 377768 439634
rect 377448 439366 377768 439398
rect 300648 435454 300968 435486
rect 300648 435218 300690 435454
rect 300926 435218 300968 435454
rect 300648 435134 300968 435218
rect 300648 434898 300690 435134
rect 300926 434898 300968 435134
rect 300648 434866 300968 434898
rect 331368 435454 331688 435486
rect 331368 435218 331410 435454
rect 331646 435218 331688 435454
rect 331368 435134 331688 435218
rect 331368 434898 331410 435134
rect 331646 434898 331688 435134
rect 331368 434866 331688 434898
rect 362088 435454 362408 435486
rect 362088 435218 362130 435454
rect 362366 435218 362408 435454
rect 362088 435134 362408 435218
rect 362088 434898 362130 435134
rect 362366 434898 362408 435134
rect 362088 434866 362408 434898
rect 285288 403954 285608 403986
rect 285288 403718 285330 403954
rect 285566 403718 285608 403954
rect 285288 403634 285608 403718
rect 285288 403398 285330 403634
rect 285566 403398 285608 403634
rect 285288 403366 285608 403398
rect 316008 403954 316328 403986
rect 316008 403718 316050 403954
rect 316286 403718 316328 403954
rect 316008 403634 316328 403718
rect 316008 403398 316050 403634
rect 316286 403398 316328 403634
rect 316008 403366 316328 403398
rect 346728 403954 347048 403986
rect 346728 403718 346770 403954
rect 347006 403718 347048 403954
rect 346728 403634 347048 403718
rect 346728 403398 346770 403634
rect 347006 403398 347048 403634
rect 346728 403366 347048 403398
rect 377448 403954 377768 403986
rect 377448 403718 377490 403954
rect 377726 403718 377768 403954
rect 377448 403634 377768 403718
rect 377448 403398 377490 403634
rect 377726 403398 377768 403634
rect 377448 403366 377768 403398
rect 300648 399454 300968 399486
rect 300648 399218 300690 399454
rect 300926 399218 300968 399454
rect 300648 399134 300968 399218
rect 300648 398898 300690 399134
rect 300926 398898 300968 399134
rect 300648 398866 300968 398898
rect 331368 399454 331688 399486
rect 331368 399218 331410 399454
rect 331646 399218 331688 399454
rect 331368 399134 331688 399218
rect 331368 398898 331410 399134
rect 331646 398898 331688 399134
rect 331368 398866 331688 398898
rect 362088 399454 362408 399486
rect 362088 399218 362130 399454
rect 362366 399218 362408 399454
rect 362088 399134 362408 399218
rect 362088 398898 362130 399134
rect 362366 398898 362408 399134
rect 362088 398866 362408 398898
rect 285288 367954 285608 367986
rect 285288 367718 285330 367954
rect 285566 367718 285608 367954
rect 285288 367634 285608 367718
rect 285288 367398 285330 367634
rect 285566 367398 285608 367634
rect 285288 367366 285608 367398
rect 316008 367954 316328 367986
rect 316008 367718 316050 367954
rect 316286 367718 316328 367954
rect 316008 367634 316328 367718
rect 316008 367398 316050 367634
rect 316286 367398 316328 367634
rect 316008 367366 316328 367398
rect 346728 367954 347048 367986
rect 346728 367718 346770 367954
rect 347006 367718 347048 367954
rect 346728 367634 347048 367718
rect 346728 367398 346770 367634
rect 347006 367398 347048 367634
rect 346728 367366 347048 367398
rect 377448 367954 377768 367986
rect 377448 367718 377490 367954
rect 377726 367718 377768 367954
rect 377448 367634 377768 367718
rect 377448 367398 377490 367634
rect 377726 367398 377768 367634
rect 377448 367366 377768 367398
rect 300648 363454 300968 363486
rect 300648 363218 300690 363454
rect 300926 363218 300968 363454
rect 300648 363134 300968 363218
rect 300648 362898 300690 363134
rect 300926 362898 300968 363134
rect 300648 362866 300968 362898
rect 331368 363454 331688 363486
rect 331368 363218 331410 363454
rect 331646 363218 331688 363454
rect 331368 363134 331688 363218
rect 331368 362898 331410 363134
rect 331646 362898 331688 363134
rect 331368 362866 331688 362898
rect 362088 363454 362408 363486
rect 362088 363218 362130 363454
rect 362366 363218 362408 363454
rect 362088 363134 362408 363218
rect 362088 362898 362130 363134
rect 362366 362898 362408 363134
rect 362088 362866 362408 362898
rect 273115 336020 273181 336021
rect 271643 333300 271709 333301
rect 271643 333236 271644 333300
rect 271708 333236 271709 333300
rect 271643 333235 271709 333236
rect 268883 326364 268949 326365
rect 268883 326300 268884 326364
rect 268948 326300 268949 326364
rect 268883 326299 268949 326300
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 232954 267914 268398
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 267294 196954 267914 232398
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 309454 272414 336000
rect 273115 335956 273116 336020
rect 273180 335956 273181 336020
rect 273115 335955 273181 335956
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 313954 276914 336000
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 241954 276914 277398
rect 276294 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 276914 241954
rect 276294 241634 276914 241718
rect 276294 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 276914 241634
rect 276294 205954 276914 241398
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 318454 281414 336000
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 210454 281414 245898
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 322954 285914 336000
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 214954 285914 250398
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 327454 290414 336000
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 331954 294914 336000
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 223954 294914 259398
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 300454 299414 336000
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 228454 299414 263898
rect 298794 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 299414 228454
rect 298794 228134 299414 228218
rect 298794 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 299414 228134
rect 298794 192454 299414 227898
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 304954 303914 336000
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 232954 303914 268398
rect 303294 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 303914 232954
rect 303294 232634 303914 232718
rect 303294 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 303914 232634
rect 303294 196954 303914 232398
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 124954 303914 160398
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 309454 308414 336000
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 313954 312914 336000
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 241954 312914 277398
rect 312294 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 312914 241954
rect 312294 241634 312914 241718
rect 312294 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 312914 241634
rect 312294 205954 312914 241398
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 169954 312914 205398
rect 312294 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 312914 169954
rect 312294 169634 312914 169718
rect 312294 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 312914 169634
rect 312294 133954 312914 169398
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 318454 317414 336000
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 210454 317414 245898
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 174454 317414 209898
rect 316794 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 317414 174454
rect 316794 174134 317414 174218
rect 316794 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 317414 174134
rect 316794 138454 317414 173898
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 322954 321914 336000
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 214954 321914 250398
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 321294 178954 321914 214398
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 142954 321914 178398
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 327454 326414 336000
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 331954 330914 336000
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 223954 330914 259398
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 187954 330914 223398
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 151954 330914 187398
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 300454 335414 336000
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 228454 335414 263898
rect 334794 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 335414 228454
rect 334794 228134 335414 228218
rect 334794 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 335414 228134
rect 334794 192454 335414 227898
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 304954 339914 336000
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 232954 339914 268398
rect 339294 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 339914 232954
rect 339294 232634 339914 232718
rect 339294 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 339914 232634
rect 339294 196954 339914 232398
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 124954 339914 160398
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 309454 344414 336000
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 313954 348914 336000
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 241954 348914 277398
rect 348294 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 348914 241954
rect 348294 241634 348914 241718
rect 348294 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 348914 241634
rect 348294 205954 348914 241398
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 318454 353414 336000
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 210454 353414 245898
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 322954 357914 336000
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 214954 357914 250398
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 327454 362414 336000
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 331954 366914 336000
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 300454 371414 336000
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 304954 375914 336000
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 309454 380414 336000
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 313954 384914 336000
rect 385174 331805 385234 457403
rect 385171 331804 385237 331805
rect 385171 331740 385172 331804
rect 385236 331740 385237 331804
rect 385171 331739 385237 331740
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 318454 389414 336000
rect 389590 330445 389650 457403
rect 392808 435454 393128 435486
rect 392808 435218 392850 435454
rect 393086 435218 393128 435454
rect 392808 435134 393128 435218
rect 392808 434898 392850 435134
rect 393086 434898 393128 435134
rect 392808 434866 393128 434898
rect 392808 399454 393128 399486
rect 392808 399218 392850 399454
rect 393086 399218 393128 399454
rect 392808 399134 393128 399218
rect 392808 398898 392850 399134
rect 393086 398898 393128 399134
rect 392808 398866 393128 398898
rect 392808 363454 393128 363486
rect 392808 363218 392850 363454
rect 393086 363218 393128 363454
rect 392808 363134 393128 363218
rect 392808 362898 392850 363134
rect 393086 362898 393128 363134
rect 392808 362866 393128 362898
rect 389587 330444 389653 330445
rect 389587 330380 389588 330444
rect 389652 330380 389653 330444
rect 389587 330379 389653 330380
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 322954 393914 336000
rect 394006 329085 394066 457403
rect 397502 337381 397562 457403
rect 397499 337380 397565 337381
rect 397499 337316 397500 337380
rect 397564 337316 397565 337380
rect 397499 337315 397565 337316
rect 394003 329084 394069 329085
rect 394003 329020 394004 329084
rect 394068 329020 394069 329084
rect 394003 329019 394069 329020
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 327454 398414 336000
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 398790 149157 398850 457403
rect 401550 338061 401610 457403
rect 401547 338060 401613 338061
rect 401547 337996 401548 338060
rect 401612 337996 401613 338060
rect 401547 337995 401613 337996
rect 402294 331954 402914 336000
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 398787 149156 398853 149157
rect 398787 149092 398788 149156
rect 398852 149092 398853 149156
rect 398787 149091 398853 149092
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 403022 96661 403082 457403
rect 403019 96660 403085 96661
rect 403019 96596 403020 96660
rect 403084 96596 403085 96660
rect 403019 96595 403085 96596
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 405782 44301 405842 457403
rect 408168 439954 408488 439986
rect 408168 439718 408210 439954
rect 408446 439718 408488 439954
rect 408168 439634 408488 439718
rect 408168 439398 408210 439634
rect 408446 439398 408488 439634
rect 408168 439366 408488 439398
rect 408168 403954 408488 403986
rect 408168 403718 408210 403954
rect 408446 403718 408488 403954
rect 408168 403634 408488 403718
rect 408168 403398 408210 403634
rect 408446 403398 408488 403634
rect 408168 403366 408488 403398
rect 408168 367954 408488 367986
rect 408168 367718 408210 367954
rect 408446 367718 408488 367954
rect 408168 367634 408488 367718
rect 408168 367398 408210 367634
rect 408446 367398 408488 367634
rect 408168 367366 408488 367398
rect 406794 300454 407414 336000
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 408726 58037 408786 457403
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 411294 304954 411914 336000
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 408723 58036 408789 58037
rect 408723 57972 408724 58036
rect 408788 57972 408789 58036
rect 408723 57971 408789 57972
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 405779 44300 405845 44301
rect 405779 44236 405780 44300
rect 405844 44236 405845 44300
rect 405779 44235 405845 44236
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 309454 416414 336000
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 118826 228218 119062 228454
rect 119146 228218 119382 228454
rect 118826 227898 119062 228134
rect 119146 227898 119382 228134
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 118826 120218 119062 120454
rect 119146 120218 119382 120454
rect 118826 119898 119062 120134
rect 119146 119898 119382 120134
rect 118826 84218 119062 84454
rect 119146 84218 119382 84454
rect 118826 83898 119062 84134
rect 119146 83898 119382 84134
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 123326 232718 123562 232954
rect 123646 232718 123882 232954
rect 123326 232398 123562 232634
rect 123646 232398 123882 232634
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 123326 124718 123562 124954
rect 123646 124718 123882 124954
rect 123326 124398 123562 124634
rect 123646 124398 123882 124634
rect 123326 88718 123562 88954
rect 123646 88718 123882 88954
rect 123326 88398 123562 88634
rect 123646 88398 123882 88634
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 132326 241718 132562 241954
rect 132646 241718 132882 241954
rect 132326 241398 132562 241634
rect 132646 241398 132882 241634
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 132326 169718 132562 169954
rect 132646 169718 132882 169954
rect 132326 169398 132562 169634
rect 132646 169398 132882 169634
rect 132326 133718 132562 133954
rect 132646 133718 132882 133954
rect 132326 133398 132562 133634
rect 132646 133398 132882 133634
rect 132326 97718 132562 97954
rect 132646 97718 132882 97954
rect 132326 97398 132562 97634
rect 132646 97398 132882 97634
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 136826 246218 137062 246454
rect 137146 246218 137382 246454
rect 136826 245898 137062 246134
rect 137146 245898 137382 246134
rect 136826 210218 137062 210454
rect 137146 210218 137382 210454
rect 136826 209898 137062 210134
rect 137146 209898 137382 210134
rect 136826 174218 137062 174454
rect 137146 174218 137382 174454
rect 136826 173898 137062 174134
rect 137146 173898 137382 174134
rect 136826 138218 137062 138454
rect 137146 138218 137382 138454
rect 136826 137898 137062 138134
rect 137146 137898 137382 138134
rect 136826 102218 137062 102454
rect 137146 102218 137382 102454
rect 136826 101898 137062 102134
rect 137146 101898 137382 102134
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 141326 214718 141562 214954
rect 141646 214718 141882 214954
rect 141326 214398 141562 214634
rect 141646 214398 141882 214634
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 141326 142718 141562 142954
rect 141646 142718 141882 142954
rect 141326 142398 141562 142634
rect 141646 142398 141882 142634
rect 141326 106718 141562 106954
rect 141646 106718 141882 106954
rect 141326 106398 141562 106634
rect 141646 106398 141882 106634
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 150326 223718 150562 223954
rect 150646 223718 150882 223954
rect 150326 223398 150562 223634
rect 150646 223398 150882 223634
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 150326 151718 150562 151954
rect 150646 151718 150882 151954
rect 150326 151398 150562 151634
rect 150646 151398 150882 151634
rect 150326 115718 150562 115954
rect 150646 115718 150882 115954
rect 150326 115398 150562 115634
rect 150646 115398 150882 115634
rect 150326 79718 150562 79954
rect 150646 79718 150882 79954
rect 150326 79398 150562 79634
rect 150646 79398 150882 79634
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 154826 228218 155062 228454
rect 155146 228218 155382 228454
rect 154826 227898 155062 228134
rect 155146 227898 155382 228134
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 154826 120218 155062 120454
rect 155146 120218 155382 120454
rect 154826 119898 155062 120134
rect 155146 119898 155382 120134
rect 154826 84218 155062 84454
rect 155146 84218 155382 84454
rect 154826 83898 155062 84134
rect 155146 83898 155382 84134
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 159326 232718 159562 232954
rect 159646 232718 159882 232954
rect 159326 232398 159562 232634
rect 159646 232398 159882 232634
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 159326 160718 159562 160954
rect 159646 160718 159882 160954
rect 159326 160398 159562 160634
rect 159646 160398 159882 160634
rect 159326 124718 159562 124954
rect 159646 124718 159882 124954
rect 159326 124398 159562 124634
rect 159646 124398 159882 124634
rect 159326 88718 159562 88954
rect 159646 88718 159882 88954
rect 159326 88398 159562 88634
rect 159646 88398 159882 88634
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 168326 241718 168562 241954
rect 168646 241718 168882 241954
rect 168326 241398 168562 241634
rect 168646 241398 168882 241634
rect 168326 205718 168562 205954
rect 168646 205718 168882 205954
rect 168326 205398 168562 205634
rect 168646 205398 168882 205634
rect 168326 169718 168562 169954
rect 168646 169718 168882 169954
rect 168326 169398 168562 169634
rect 168646 169398 168882 169634
rect 168326 133718 168562 133954
rect 168646 133718 168882 133954
rect 168326 133398 168562 133634
rect 168646 133398 168882 133634
rect 168326 97718 168562 97954
rect 168646 97718 168882 97954
rect 168326 97398 168562 97634
rect 168646 97398 168882 97634
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 172826 246218 173062 246454
rect 173146 246218 173382 246454
rect 172826 245898 173062 246134
rect 173146 245898 173382 246134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 172826 138218 173062 138454
rect 173146 138218 173382 138454
rect 172826 137898 173062 138134
rect 173146 137898 173382 138134
rect 172826 102218 173062 102454
rect 173146 102218 173382 102454
rect 172826 101898 173062 102134
rect 173146 101898 173382 102134
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 177326 106718 177562 106954
rect 177646 106718 177882 106954
rect 177326 106398 177562 106634
rect 177646 106398 177882 106634
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 190826 228218 191062 228454
rect 191146 228218 191382 228454
rect 190826 227898 191062 228134
rect 191146 227898 191382 228134
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 239250 435218 239486 435454
rect 239250 434898 239486 435134
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 239250 399218 239486 399454
rect 239250 398898 239486 399134
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 239250 363218 239486 363454
rect 239250 362898 239486 363134
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 231326 232718 231562 232954
rect 231646 232718 231882 232954
rect 231326 232398 231562 232634
rect 231646 232398 231882 232634
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 240326 241718 240562 241954
rect 240646 241718 240882 241954
rect 240326 241398 240562 241634
rect 240646 241398 240882 241634
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 254610 439718 254846 439954
rect 254610 439398 254846 439634
rect 254610 403718 254846 403954
rect 254610 403398 254846 403634
rect 254610 367718 254846 367954
rect 254610 367398 254846 367634
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 269970 435218 270206 435454
rect 269970 434898 270206 435134
rect 269970 399218 270206 399454
rect 269970 398898 270206 399134
rect 269970 363218 270206 363454
rect 269970 362898 270206 363134
rect 285330 439718 285566 439954
rect 285330 439398 285566 439634
rect 316050 439718 316286 439954
rect 316050 439398 316286 439634
rect 346770 439718 347006 439954
rect 346770 439398 347006 439634
rect 377490 439718 377726 439954
rect 377490 439398 377726 439634
rect 300690 435218 300926 435454
rect 300690 434898 300926 435134
rect 331410 435218 331646 435454
rect 331410 434898 331646 435134
rect 362130 435218 362366 435454
rect 362130 434898 362366 435134
rect 285330 403718 285566 403954
rect 285330 403398 285566 403634
rect 316050 403718 316286 403954
rect 316050 403398 316286 403634
rect 346770 403718 347006 403954
rect 346770 403398 347006 403634
rect 377490 403718 377726 403954
rect 377490 403398 377726 403634
rect 300690 399218 300926 399454
rect 300690 398898 300926 399134
rect 331410 399218 331646 399454
rect 331410 398898 331646 399134
rect 362130 399218 362366 399454
rect 362130 398898 362366 399134
rect 285330 367718 285566 367954
rect 285330 367398 285566 367634
rect 316050 367718 316286 367954
rect 316050 367398 316286 367634
rect 346770 367718 347006 367954
rect 346770 367398 347006 367634
rect 377490 367718 377726 367954
rect 377490 367398 377726 367634
rect 300690 363218 300926 363454
rect 300690 362898 300926 363134
rect 331410 363218 331646 363454
rect 331410 362898 331646 363134
rect 362130 363218 362366 363454
rect 362130 362898 362366 363134
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 276326 241718 276562 241954
rect 276646 241718 276882 241954
rect 276326 241398 276562 241634
rect 276646 241398 276882 241634
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 298826 228218 299062 228454
rect 299146 228218 299382 228454
rect 298826 227898 299062 228134
rect 299146 227898 299382 228134
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 303326 232718 303562 232954
rect 303646 232718 303882 232954
rect 303326 232398 303562 232634
rect 303646 232398 303882 232634
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 312326 241718 312562 241954
rect 312646 241718 312882 241954
rect 312326 241398 312562 241634
rect 312646 241398 312882 241634
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 312326 169718 312562 169954
rect 312646 169718 312882 169954
rect 312326 169398 312562 169634
rect 312646 169398 312882 169634
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 316826 174218 317062 174454
rect 317146 174218 317382 174454
rect 316826 173898 317062 174134
rect 317146 173898 317382 174134
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 334826 228218 335062 228454
rect 335146 228218 335382 228454
rect 334826 227898 335062 228134
rect 335146 227898 335382 228134
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 339326 232718 339562 232954
rect 339646 232718 339882 232954
rect 339326 232398 339562 232634
rect 339646 232398 339882 232634
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 348326 241718 348562 241954
rect 348646 241718 348882 241954
rect 348326 241398 348562 241634
rect 348646 241398 348882 241634
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 392850 435218 393086 435454
rect 392850 434898 393086 435134
rect 392850 399218 393086 399454
rect 392850 398898 393086 399134
rect 392850 363218 393086 363454
rect 392850 362898 393086 363134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 408210 439718 408446 439954
rect 408210 439398 408446 439634
rect 408210 403718 408446 403954
rect 408210 403398 408446 403634
rect 408210 367718 408446 367954
rect 408210 367398 408446 367634
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 254610 439954
rect 254846 439718 285330 439954
rect 285566 439718 316050 439954
rect 316286 439718 346770 439954
rect 347006 439718 377490 439954
rect 377726 439718 408210 439954
rect 408446 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 254610 439634
rect 254846 439398 285330 439634
rect 285566 439398 316050 439634
rect 316286 439398 346770 439634
rect 347006 439398 377490 439634
rect 377726 439398 408210 439634
rect 408446 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 239250 435454
rect 239486 435218 269970 435454
rect 270206 435218 300690 435454
rect 300926 435218 331410 435454
rect 331646 435218 362130 435454
rect 362366 435218 392850 435454
rect 393086 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 239250 435134
rect 239486 434898 269970 435134
rect 270206 434898 300690 435134
rect 300926 434898 331410 435134
rect 331646 434898 362130 435134
rect 362366 434898 392850 435134
rect 393086 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 254610 403954
rect 254846 403718 285330 403954
rect 285566 403718 316050 403954
rect 316286 403718 346770 403954
rect 347006 403718 377490 403954
rect 377726 403718 408210 403954
rect 408446 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 254610 403634
rect 254846 403398 285330 403634
rect 285566 403398 316050 403634
rect 316286 403398 346770 403634
rect 347006 403398 377490 403634
rect 377726 403398 408210 403634
rect 408446 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 239250 399454
rect 239486 399218 269970 399454
rect 270206 399218 300690 399454
rect 300926 399218 331410 399454
rect 331646 399218 362130 399454
rect 362366 399218 392850 399454
rect 393086 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 239250 399134
rect 239486 398898 269970 399134
rect 270206 398898 300690 399134
rect 300926 398898 331410 399134
rect 331646 398898 362130 399134
rect 362366 398898 392850 399134
rect 393086 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 254610 367954
rect 254846 367718 285330 367954
rect 285566 367718 316050 367954
rect 316286 367718 346770 367954
rect 347006 367718 377490 367954
rect 377726 367718 408210 367954
rect 408446 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 254610 367634
rect 254846 367398 285330 367634
rect 285566 367398 316050 367634
rect 316286 367398 346770 367634
rect 347006 367398 377490 367634
rect 377726 367398 408210 367634
rect 408446 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 239250 363454
rect 239486 363218 269970 363454
rect 270206 363218 300690 363454
rect 300926 363218 331410 363454
rect 331646 363218 362130 363454
rect 362366 363218 392850 363454
rect 393086 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 239250 363134
rect 239486 362898 269970 363134
rect 270206 362898 300690 363134
rect 300926 362898 331410 363134
rect 331646 362898 362130 363134
rect 362366 362898 392850 363134
rect 393086 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use user_proj_example  mprj
timestamp 0
transform 1 0 235000 0 1 338000
box 1066 0 178886 120000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 336000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 460000 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 336000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 460000 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 336000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 460000 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 336000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 460000 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 336000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 460000 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 336000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 460000 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 336000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 460000 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 336000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 460000 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 336000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 460000 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 336000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 460000 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 336000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 460000 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 336000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 460000 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 336000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 460000 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 336000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 460000 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 336000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 460000 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 336000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 460000 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 336000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 460000 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 336000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 460000 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 336000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 460000 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 336000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 460000 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 336000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 460000 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 336000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 460000 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 336000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 460000 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 336000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 460000 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 336000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 460000 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 336000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 460000 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 336000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 460000 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 336000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 460000 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 336000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 460000 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 336000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 460000 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 336000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 460000 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 336000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 460000 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 336000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 460000 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 336000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 460000 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 336000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 460000 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 336000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 460000 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 336000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 460000 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 336000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 460000 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 336000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 460000 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 336000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 460000 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 336000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 460000 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
